LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.std_logic_textio.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

LIBRARY STD;
USE STD.textio.all;

entity Decoder_TB is
end entity;

architecture Decoder_TB_arch of Decoder_TB is

component Decoder is
		port(  
		clock  : in std_logic;
		input  : std_logic_vector(254 downto 0);
		output : out std_logic_vector(254 downto 0)
		);
end component;

--TB clock
signal Clock, ok : std_logic;
constant clk_period: time:=10 ns;
signal result : std_logic_vector(254 downto 0);
signal test, check  : std_logic_vector(254 downto 0);
signal counter : integer range 1 to 4;

--FOR SINGLE TESTING
--type ROM_type is array (0 to 0) of std_logic_vector(254 downto 0);
--constant ROM_R : ROM_type := ( 
--0 =>  "001010000011101101110101001010011110001010111010110011010011001111000111110001110010010001100010011101100010111011001011111110011010001011100101111101110010010001000001110010000010101100100000101100011100111001001010010110110101101011110100101001100100000"
--);
--constant ROM_C : ROM_type := ( 
--0 => "001010000011101101110101001010011110001010111010110011010011001111000111110001110010010001100010011101100010111011001011111110011010001011100101111101110010010001000001110010000010101100100000101100111100111001001010010110110101101010110100101001100100000"
--);


type ROM_type is array (1 to 4) of std_logic_vector(254 downto 0);

constant ROM_C : ROM_type := ( --REVERSE(C)
1 => "010111001111110111110010011101111001110011100010101011100000001001101110010101000010111111110000100101010001110111010100010001001010000111100010001100011100011010000011110101111001100001111011110010100111000110111100100000001101011100011100111001010101100",
2 => "011101100101101100000011111010111100011111110001111100010000110010101101101110011010011101100110101000000111000000010100000010111110001000000111010110000011011001111001101100100101011000101110100111011000111010001011111100011100100100110001001111100001110",
3 => "111011010001011010110011101110111010111001101101110001110001011100110010011010100101111100010111001000100010011101010110100001110100011110101111101000111101010011000101110000110010011011101010010001111100110011101100101011101011110111001011111100000001100",
4 => "101100111101001101000110000001110000001000001110000001011011111110001011111110000000011110010011010001000011110100101001100110010110000001101101000011010000011100010101101010010001010110101111101001101000101001100111010101110100000000111100100011101100111"
);

constant ROM_R : ROM_type := ( --REVERSE(R)
1 => "010111001111110111110000011101111001110011100010101011100000001001101110010101000010111111110000100101010001110111010100010001001010000111100010001100011100011010001011110101111001100001111011110010100111000110111100100000001101011100011100111001010101100",
2 => "011101100101101100000011111010111100011111110001111100010000110010101101101110011010011101100110101000000111000000010100000010111110001000000111010110000011011001111001101100100101011000101110100111011000111010001011111000011110100100110001001111100001110",
3 => "111011010001011010110001101110111010111001101001110001110001011100110010011010100101111100010111001000100010011101010110100001110100011110101111101000111101010011000101110000110010011011101010010001111100110011101100101011101011110111001011111100000001100",
4 => "101100111101001101000110000011110000001000001110000001011011111110001011111110000000011110010011010001000011110100101001100100010110000001101101000011010000011100010101101010010001010110101111101001101000101001100111010101110100000000111100100011101100111"
);


begin

CLOCK_PROGRESS : process
	begin
		Clock<='0';
		wait for clk_period/2;
		Clock<='1';
		wait for clk_period/2;
end process;

tester : process (Clock)
begin

	--test <= ROM_R(0);
	--check <= ROM_C(0);

	if (counter = 4) then
		counter <= 1;
		test <= ROM_R(counter);
		check <= ROM_C(counter);
	else
		counter <= counter + 1;
		test <= ROM_R(counter);
		check <= ROM_C(counter);
	end if;

end process;


checker : process (Clock,result)
begin
	if (result = check) then
		ok <= '1';
	else
		ok <= '0';
	end if;
end process;


dut : Decoder
	port map(
		clock  => Clock,
		input	=> test,
		output => result
	);

end architecture;

