LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.std_logic_textio.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

LIBRARY STD;
USE STD.textio.all;

entity Decoder_TB is
end entity;

architecture Decoder_TB_arch of Decoder_TB is

component Decoder is
		port(  
		clock  : in std_logic;
		input  : std_logic_vector(254 downto 0);
		output : out std_logic_vector(254 downto 0)
		);
end component;

--TB clock
signal Clock, ok : std_logic;
constant clk_period: time:=10 ns;
signal result : std_logic_vector(254 downto 0);
signal test, check  : std_logic_vector(254 downto 0);
signal counter : integer range 1 to 100;

--FOR SINGLE TESTING
--type ROM_type is array (0 to 0) of std_logic_vector(254 downto 0);
--constant ROM_R : ROM_type := ( 
--0 =>  "001010000011101101110101001010011110001010111010110011010011001111000111110001110010010001100010011101100010111011001011111110011010001011100101111101110010010001000001110010000010101100100000101100011100111001001010010110110101101011110100101001100100000"
--);
--constant ROM_C : ROM_type := ( 
--0 => "001010000011101101110101001010011110001010111010110011010011001111000111110001110010010001100010011101100010111011001011111110011010001011100101111101110010010001000001110010000010101100100000101100111100111001001010010110110101101010110100101001100100000"
--);


type ROM_type is array (1 to 100) of std_logic_vector(254 downto 0);
constant ROM_C : ROM_type := ( 1 => "010000101010111001010100011011110000010111110110110010111111001111110111110001000100110111101011101100010110111111001001111101000101011101000101100111001011011011110111110100111101101101111101010011111111010110011101000100100000010011100010110010011111101",
2 => "110110011110111100000010110001111101111111001001101001010001011011000010110010010101000001000001111001110100101011001100011111010010011010101110101011010101000110110110010111110001111001011001101111110010111111111101000101100011110010111001011000100111110",
3 => "111000011110011110000000001100110011000110101010000010100010110010101101011100101110101111111001101010011011101011100001100000010101001101001101000001110110101110100110001100101111110010011000101001110010101111011001101000000000000101100110100111111100110",
4 => "011111100011011100001011100001011101011111000100101111101111111010011100010000111111000000011010100000101100000101101011111000100111000000010110011011100010011100011100011101001001101011101111010010100101100001000011110000111110100100001111111101001100010",
5 => "111011100000111011011101110111000001011101001110001111010111100110111110111011000010111100100010101010101010100100101001111100111001101001101001001000011000000001110010011101011110011000001001111010010000001111000101001111010110110010100001001101010100001",
6 => "101111101001100110100011100001011110010000110010100010000100100110010000000001011011011010011011000000011011000001000101001000111111001000101110101010101110000100010101000000011110111101010000100001000010011010110100010000101101000000101000100010101101101",
7 => "010110110101110101011000001101001010001110100011011001001101111010110000100110011011111101110100001001101110111000011011111100111010011000110111011010100010000011101111110001000000111110010001111100000100011000011101100010111110101000101001110011111110010",
8 => "011111011000111111100011101000011000111100101101110011011100010011110001110011001100101010010000111111101100000000100110101100110000110000000100000100010010100011100001111111011100001111110110110011011000101011010001100110000000010010111101001011000000010",
9 => "101111011011010000101111010111101110101000101111111010111101011100001100101010100010010000111111110001001000000100111111010011111011000110010000011001111100111000111111001011111011100101100010101111100001100000011110001111100001011000111010100111110010110",
10 => "101011011111011010111101010000111110000000101101100011011000000010000101010100110101001000011110001100000101100110100011001111011001111010001111111001001000110111001001101011010110111001111011001000101011010101011000100100011000000011010011000010000101101",
11 => "101110110011011000010011000000000100001010001010101101111111001011111000111000101001101110111000111111000111000000001010000111111100100000111000101101110010101100001110100111000100011010111011001110010101000010011101011100011001101011110011011100001000100",
12 => "110000110101000010001011000001011010110110000101001010010101000010000000010100011010101100101010010111000011000111010001010101011010010110000100010001011000111110000101110111000101001101100110001101110101010111100111100111001111011010111000101010010111101",
13 => "010000011011110101101100110100110110100000101001101000010000011101000100000101101101101010100001101010011001011111000100111001101000001000110101000001101011111000111000010010100011110001011111011110010000011111101110100011011101110101000001000100110000010",
14 => "100111001100010000010011100110001100000001111111010001010111000100110110000001110001110011101000110001111111101111110001111001101001100000001011100100111100101101100100101010011110110101010100101101110100001011010010110110100100000111110101000101110000101",
15 => "101111100100111011111111101111101110101110101001101001111111001010111000101100111110111101010101010011010100100000111110101010110001101101111111000000101111010110001101110010101000100111111001001000000100110110101000000011000110110111100101101011111011001",
16 => "000000100010101010101010111101100000001010001110011011110000000100000100111001100000001111001100010011110001100100111000111111101110110001110111000010111110001100101100110011011000000001010001001010000110001111100011110100011100011001001000100100101010011",
17 => "101001110010111011110111100001110101011111111111101100111000010001110100110001101000100100000001011101110011000011011000000100100110001110011100001010111000110110010110110100111101010001010011111110101010111010111111011100001110101010100100011100000010011",
18 => "111110101100111001100101111100110011001110000110001011000010010011010001011101110110110100011101100011101000011111110011011101010110110011011011001010101011010111110101101101101100000011010000001010011100010010001000000111000000001110101110001011000110110",
19 => "001111111101010000000101001100000011110110100000000000011011001101100100111001001111111111010110001111110100111100101010011101000001001100100000011000111101010011001001010001100110111101101011010100110001010001011110011110011101110000101010011100101101010",
20 => "100010000001101001101000111100101111010000010001010011101000011100111001100100111010101000010001110101111001101100000110000100101001111000000001001110111001110111000100000000110100100110100111001011011101111001111100000100100111101111000010001111110001011",
21 => "111010010111101100111111101110101000100011111100011110111000101000101100010001010001010000111001100010111111000100000010101011111011111001010110001000000101111101110000000101011100101111111101001010101111100111110010001110000000001000011010100000001110011",
22 => "000100010100000010100111101011111110011110000100000111100101011000011111110101100000001111011010101111001011000111101101111000110110011010100101010011101101010001001010001001110001111111101101011100110000111111000001111100100000001111000001110111010000011",
23 => "110000010111001111111100101000111011101000110000110111000110110000101011111111111000000000101111100101100110000001100100111011101111101110011101111000011000100111110111100011000011010100001011010000011010001111100101001100010000101111010110011000001011010",
24 => "111110000000011001011000111010000100111110010001101111011001000101001110000010100110001100110000010011111111111111110010101000111001101111010001000001111001010101001011001111100000110110000000101010011010001100001000000101101101011110111011100001000010100",
25 => "111101111111000100000010100110101000110101101001010111001010111000001010011100000101111010101010000111110010100110011010100010111001100100101001001111011111010100100100011010100001011011110110001010111111000010111000100110000100001011111000101101011010000",
26 => "100010100000001110011000110010010111011101110100110100100011111001011100000011101001011011101110110001001010010111110100100010001111000101010001001010010010000011010110111001110111100100100110011001000010110000011001110100100110111001011101001000101000010",
27 => "110001110000001011000101101111001100110101010010011100101100110100110001110010110111001010010011111110110110100011000001010010100011111111010110101010100011100111101110100101000101100110111101101110110100111010011011010001111111010101110111111000100001110",
28 => "001001010011000011010000101100001111001011100001000010100001101011111100100000010101110111110011001000100101010010000011110011011101111101010110001101000001111100101111011001001111110010000001101001011001001100001110010000010010100101100101011001101111111",
29 => "001011100011011101001101010011110010011001111010001100101110011111100010101000111010101010100100111101010111000011101000001101101010100100101011001001100000111001111001111100001010101111010011000110110100111111010000011110110010101100110011111011011110001",
30 => "011010011001110010000011000101100110101101011100101111100111010101000011000101001110100000000100111101000100010111011000101110000100010001110101010101011110111001011000100100111100010110010001010101010100101110010010001011111100001100011111001010100101110",
31 => "010101111111000010000101111001110111011110101001000011111001101110111001101011011101011100100100010010111100001001010011111111101000100100111111100011111001110001011101010111100010000101111101011000110100111010110111100001110001010100100000100101001010001",
32 => "110010100110010111111101000010000000001000000111100011010000111101010110111101000011001101000000010000010111001110010001001101101010011011100101110110100111011101010101100101101101000100101101001101011001100001111101110011001011111010001010000011110100001",
33 => "111010101100101110001010011101100100101000000100000001110110101011111100001101110101111100001001011000000001011000001111010011110110101110010111101001110110111011101010100110100111011110111000010011111001001110101000001110101011110011010001100010110110010",
34 => "011110111001110110101100101000010000001101110100001001010010000101001110000101000010000000011101011011000111101110000111100001000000111101101111001110110011011110110011101011001101010010000001010001101011001111111100111010011011110011111110011101001011000",
35 => "100101001010101001001101011111101011001000001000101100010010110010101001100110100000000000110011010100100101010000111111001111100101101011100000101011110100101001011101001100110110110110100100111111000100001111101011000000101101010010001010101011001010110",
36 => "001100011011000111101010000010001010001011110000100000100110010100111011000011111010010010110100111100001010111011001100110000100000000001100010010101001010100111100000001010111001101000100110000101001011001101100100001101000110000010110001001011111111101",
37 => "100001111101011110000010111011011011011000100101011100010111000101100100100100100101100110000110101101111010010000001000101011000000100111100010101100111110111000100111010110110100001111111001001101100100000000001100001010111010100001010101110100101101010",
38 => "100000011101010001011110101001001101000101000010001001011001000010110001100001100101000011111011010110010101001000110101000101100001010101001010011010111001100100110010100000101000100000111011000001110011011010000010000000100111011110001010000111110001011",
39 => "100101001011010100101000111110001110011111001011111011100011011100101011100100111111101000111001100101101001010011010111001011111100001110100011000100010001111100011000110100101010010000001011111110011100000010011011111110111011000100100010100000111110010",
40 => "111101100110011011100111011000100100000100101111000001010000000101001000101110111110000100001011000111010100111001001010101110101000101110110111001100010110110000011011001100000111001000001001011111110000100001011111000010101111110000000011100111011111001",
41 => "001010100100101000001100000111111101000011011001000011111000010100010010000000100001011111011111111101011101100010010101000101010010111110001001011010101011111011000000111100101110100010011001101101011011000000011000101110100101111100100110101000100000000",
42 => "010100010110101011001100001101010010001111010000110110010101110010101010011010010111000001001100010110110101111101100010001110001011101101101101110111011000000001110101001011011100100111100001110001000100110010000110011010110010100010111011111101001001100",
43 => "111100100111100110110101110000001101100110011001100110101111110111101000100111111001010100010001110011000101000000010001001110101111000011110001100010111000111111111001010010100000011110100010001010111001001100111000001100110010101100101010110011110010111",
44 => "000000000000110010100111011001001100101110100001111100110110010101011111010010010110010101000100000011001001101011000100111101100111010010110101010101011111001111010010010001011101110100010100001011010110010110001110110011010100001011010101010011110000001",
45 => "100110001000111100010100110111011110101010000111100100101011111101101110101000000000000010001011101010011001000101001011010100100001000000011100011111100011010100101101001000111001111101011011001110100101000010011111000010110101110000010100100111001001111",
46 => "110100010101010000110111000100100101110010000011111001111010010011101111100111010000000101111001000001000011111001010110001011111010101001100001110100011001100001100101110101101111001101100011111010000000110101111101001101100001000110100001010101011101100",
47 => "110011011110111000001111011001001101000111100010011100000100000010110101101101100000100010010100100000011001101000011100010011110101010001110110100110010111000111101000010101110010110110100010011000100001011111001001001000001010000000110101110010101110010",
48 => "001010110100011000000011010101110110100101100111101110100111000110000010000100011000110010010110001111011010001010000101001010000110100101100010000011011010010101100000011010010001101000110011001110101001111100001011111000110000000011100101110111000000001",
49 => "110000000000001111000011111110011111110110111110110000010100110101110110001111110100001110101101111000110010000010010011000111100000010001001001010100011010110101000010111101011011100110100011010011110110000000010100110101101010101000011000001111100010111",
50 => "110010111111001101111001010111100100001011010001010011110110110011011110110001101010010001011100000111110101011100110101100100010101001010001101101110100111001101011101001100111111111000000100001000010010100111010000101100001100100010011010010010101011001",
51 => "111010101010110000011011111000001001010011111011010111101100111100011011010011100001110011011100110011110101110011001001001000111011110011100000001100101001000000001001011000101100011000100110100100010001110101001010110001110011100100011100110001011110100",
52 => "000000011011101111101001001111100100110110010110010101111010001111011010111101110100111010000111100011011010111111101100000111011011000111101101101001010000011100001011010101101010000001000000011111010100100101100011010111100000100110101100010110001100010",
53 => "110010110001010010010100010101110110011011111101110001111111011011100101111011101100100110110100010100101101001011110100001111001100111011100010100010110111101000110110011000101000111011111001100011111001001110110010011001000110001000101101011011110001111",
54 => "000111011101000011100100101000010001001010100011101000000010100111100000000011000110111011010010001110000011101000110011100000000001100000001010111011011110000111000111111001010100001000100011101011011010000000101000011111010011100001001011111100101100111",
55 => "101000000000011011111100110001111100111001000100011000111000100100101100110000101011111000100011000011101011101011011011101100010011000111111111101111111111001100010101011100101101010110010001010111011101100010000000010110101011111101100010100101000101100",
56 => "110010001001101010111101000001000011100010000010100110000000010011000011010001001011010011101000110000101010111010101000010101111110101111001011011110001111001110101010000101110101001010111111011000100001001111100110111111000001101000000110000110011110000",
57 => "010010111001010010100010101000101001011110011100001011101111100001111100111101110010110001101101011010011001000111100010101001101111101001000100011100000111001000110000000100000100101010000100101101011100100110011010001100110110010101101111110001010010001",
58 => "101001000110101011011011001100110010011111111001100100101011010010000000011101100001101110000101111111101010100111100101000001000010001100010001101001100010111001000110111110100011110111000111111101000010111101010000010101000010100110001111100010101101100",
59 => "111111000011101000111111001101010011101100101010111000110001001011010000001000110010101010101001010010100100110110101000101110110111110010100000111111110000000110000110000110110110011111001111010101000001111111100111100101000010101001001001011101111101111",
60 => "010110101100111000101110111001111011011110111111011101000101101010010000010001010010011000110110010100111101110111101010010011000110110000111111001100010100110111100001110111001100101100010101110110001010001010010100010111111000000100001111111000100001001",
61 => "111111000101100100010010101000111001101011001010111110001100100101011111000101111000010011010011000001010001101100110001100011010110000011111111110101100100100010011001111111111101000001000110011011010010100111010110000100111000010001011000101100000001010",
62 => "110001010000111000100111110111111000010100101110111111001000110000001000101111001110011100110010111100010100001111011001101011101101110111101010011011000100111001000101000011101001010001111101010001101100011000110100001010110001110110010000001100101010100",
63 => "011100101011010001111000101001001111000011110100010001101000010110010100110111001000110001100011101000011111000010010011010110000001000111101100011010111101001110011010001111110101111001110111100010100110011110000010011111001010000110011010111000010010011",
64 => "001001001110111000111010101110010101000111110011110000110110111001100010101100101011010111001100010101011011101001101001000111110000101101010001001000101110110110110111110110010000010011101001011111001001000000110101100110000001110110010101111011000110101",
65 => "001010101101001001100000110111110111001010011010111111101101100110011101110010011010011100100110001111011110010000010001001011110010100001110110001110011011011001001010001000001010011011101100111110110101101000101011111001100101001001110101010111101000000",
66 => "101111111000110010101111101000101100100001111111011100011101000101111110100101110110110110110111001010100010111011000001100110011111010001000011010111111100010000111010000101010101010011111100011111100101010011100100111010001000010010001110011000001011101",
67 => "101111100010001011001001000001111000111111110100011011100010101011111011101000100000000111100110011010101111010001001011000001001110100110001110010000100001101001011111000001100010101010110111101010000101111011010101101101011000110101111011000111111011000",
68 => "111001111001010011001011110010110100001000110000000101001100011011011001011111000100110010000101011111111010100100100000110011010011101100111111001011000101001100100000100011000110101101000100001000010000000000001100011110011001010001110101001001100111101",
69 => "010001011101000011000100001011011110111001101110001001010110101010111001001110110111001101100000110001100010010001010111101110000101110100111001101110000000010101101001010011011001011111110110111010011010011100001000111101000101110001010011100010001011001",
70 => "111100110110010101000010100100000010000111011010101000001100100010011101110100100101110110110101101110000010111101111111011111000110000100101011010010110001011101101100100010001010000101000100101100010100100101110010010100011000101101011100101100010100010",
71 => "011100011101010000101011010111111011100111111101010110011011100000010110000100111011110111111010000010101110111001010111100010110000001000001111001011010011000010010011100011110101001001010111001100101111010000010111010111100011011000000011100110001011111",
72 => "000010111101010101001011001100001101010111010101000001000010111011010001111110010000110110011011000000000101110000001110111011101010110110000010111001101111101110001110010011111110011011000100111010110001010001000100011111111101010010000010110101000101100",
73 => "000010010111011011001011001111000010111100111100111011010011100110110100100110111010100100011110110011111000100110101001000101110110101010001100001111011000101010000100011001111111010111011000111010000001010101010110100000100010100011000111000010010001011",
74 => "101011010101001111111011110011000000011100111010100111101111101110010101001100101100001101010001111111001010010001110000001111110001100100110100000111000101101111000001110101011011001010100010011010101110000011011010100001101101001101110101010001110110101",
75 => "100110101011100100111011011001110001101001001011001100000011110111001101010110111010101011011110101011100000011011001101100100000101111010000110011010111001101000111111100111000110010010110010001110100110010011001000100010110100101001111010111110100101011",
76 => "011101101000001010010011110001010011011100001011100000101000011000000000001001111101100101101010010001010111111010101001010001111111000101010111111100101000000010001110010011001110110100000100101011000000110001100110110011100010100110000011111101111101111",
77 => "111101110100001010101101011010111000001110100110010000010111010111000101100101101011100100010100001001010101110101001101000000000000111110100111001011001101011001101100100011110101001100000100100001101000011100111011110011011100000110010101100000110011110",
78 => "100111000010111100110000010001111000111100110111001101111100001001111111110110011010100010010010010001100001110011000100000001011010001101110111111000000000110111111101010101101101010110111011000110001010111000011101100000101110000011100010011011010001100",
79 => "001010111101011001100001101011000110001001110010110011000101011110110100110111011110101100110010011101011001010100010110100000110000010000010101101000000111110010100010110110011101110010110011001001011000000110011110000010011010110000100010110010000111010",
80 => "110111101111000100011111001111100100000011111000010001101101100001000100000100001100001011100100000111111010010111101100001101101010101101001001010001110011010001100110011010000010100101001010010001111010101110000000011011001110011100111010000110111001001",
81 => "011001011110000000111111111101101111101011110011000010101101100010011110010100101100110011001110001111100101111011010000111000101100101000110001111111000111010000111110111110001110100110011000001011110111111011111101110101011100101011100010101010100011010",
82 => "000110001101111110100101100101101110100000110101101000010101110100110000010111110000110000100110000010010111111100110010100111011011111001101110100100111010011101010111100110011000100100010000000000111010110011111111110001100010110110111001000110001001111",
83 => "001111110111101100001100101011001010010100111010111101001111010111100011011111111110111101110100010100001001011011000011100011101101111110001010001111010110000000100100100011111100000101011100111011111010001001010011001100001110100111010001011110000000110",
84 => "001110011011001010111010101001101010110000110000011001110110111111001110110101000001101101010111110001111000100100111110111001110111010111110100011110011111100010000010101010010111101011000001100010010011100010111001010000110000010010101001011110000100011",
85 => "001101101010000100101011101111011011000000110010001011101101010111111110000010011000001011001111011001100011100011011110101101011001001100111001111011000011001011101011110110111001011001011101101100011101110110110001010101100001101110001001101001110011010",
86 => "100010000000000100110001101010100110001101110001011111101010111111110000000100000010100010001111010001101100111001110001001001010001111011110001000010000110011001110011110111010101001100110100010100011110010110110101001100001011111100010011001111100001100",
87 => "110010010110010001011010000001110111100101111000000010110111011100010011011101101101000000010110000110110100101011111011101111101010100000001011101100010110001000011110000101110011011011010000001111011000010010111111001011011101010001101001101001010110101",
88 => "101111110000000111111000110100011101001110110001100001111010110011111011100110011110011001110001101011111111111010100000010111000000000110001000111111100101010101010010000011101110001011000101011110101000110001010011000110001000100110010110101100111110011",
89 => "011001010011101101110011001010100100101010101100011101000010010110111010110011110110100011100011100010100101001110101101111011110100001010101000111101011100101011001001110111010101010011111101100010110100110101011011100011000100001100001011101110011000011",
90 => "001010011100001100100110110001111101100111010111100101001010111110111001100111010100010001111010010001111000101110011110100011011001100100100100001000001100100101011110101110001000011110101111110100001100010010000001110010000110110111000001110010101100110",
91 => "111010101010010011001111011010011100011010100110101000100100011000001101000111101001100110110001101101000100101011101110000011101100011001010001100100000011000000101010111101101101100110111100011001011100110111110110101000100111110111101011001101110101001",
92 => "100110010011110001011000101100100001100000011100100100111000110101110101001100010100001111110001010011110110110001100011101001110110110000101001011001101000110010001111010010001000110001000110000000110111010011011001000011001001000000001111100001000001001",
93 => "011000110010011111101100101011000001011000110110100001011000001001001110101100001110001111110011110111001101111011101111110000101010001000100111111010001010010111010011011011111000011000111000110101000101000100011101010101101111101010010100110001001011100",
94 => "011011100110101101010110011001101101101010001111100110111010101111010010011100001100001110100010110001101010001011000010000100101010101010000001000101001000001110010011110111011110111000110010001000101010001001100000110010001111100010110010101011010010101",
95 => "010001001001001010111000011101010110111001001001001111110110101010011010110000100010001100101100000011000111100111100101110011001000111110010100101111010011010110001100000110111110010111111111110101000100110101110100101100000111111000100011000110001100100",
96 => "011011000000110011001110011010011100010101001101101101000011110011111110001110110101010100011110111011010000010111000101110101100010010110011001111111111010011000111111000110001101001011110011000101011001011001100001000001100101001101111110001001101101101",
97 => "001011110100000011100110101101000100010111001010011010101101110110011011001001110011110000110100011100111000010110010001001001011101111001101100011110100110000100110111011011011100000001000100010001100011111001001100111110110011111011000111000001100111110",
98 => "010000010111110001010100000011101011011010100001010010110000101111101000010010101000000101010011001111100011000101011001010010111010000000100011010100001010100001101110001111011000111110100100001100110111001110011010000100101110000111001010110000110000010",
99 => "011011000000100001010110011011010001100011011101111111010111101110110100011001011101000100010111010011100011110110001101000011111011001001010001011100010011111000001101110001110011001001111111011000101111010011011110010011001000111001110001010001010001100",
100 => "001001101010011011001111011011001000100000001001110100011000101001001100010011110000101100100010001010110001111100000010001111101011100110001111000001110010001111000000100100110010100011101100111000000011101101010100011011001111000000100000111101110111111"
);


constant ROM_R : ROM_type := ( 1 => "010000101010111001010100011011110000010111110110110010111111001111110111110001000000110111101011101100010110111111001001111101000101011101000101100111001011011011110111110100111101101100111101010011111111010110011101000100100000010011100010110010011111101",
2 => "110110011110111100000010110001111101111111001001101001010001011011000010010010010101000001000001111001110100101011001100011111010010011010100110101011010101000110110110010111110001111001011001101111110010111111111101000101100011110010111001011000100111110",
3 => "111000011110011110000000001100110011000110101010000010100010110010101101011100101110101111111001101010011011101011100001100000010101001101001101000001010110101110100110001100101111110010011000101011110010101111011001101000000000000101100110100111111100110",
4 => "011111100011011100001011100001011101011111000100101111101111111010011100010000111111000000011010100000101100000101101011111001100111000000010110011011100010011100011100011101001001101011101111010010100101100001000011110000111110100100001111110101001100010",
5 => "111011100000111011011101110111000001011101001110001111010111100110111110111011000000111100100010101010101010100100101001111100111001101001101001001000011000000001110010011101011110011000001000111010010000001111000101001111010110110010100001001101010100001",
6 => "101111101001100110100011100001011110010000110010100010000100100110010000000001011011011010011011000000011011000001000101001000111111001000101110101010101110000100010101000000011110111101011000100001000010011010110100010000101101000000101000100000101101101",
7 => "010110110101110101011000001101001010001110100011011001001101111010110000100110011011111101110100001101101110111000011011111100111010011000110111011010100010000011101111110001000000111110010001111100000100011000011101100010111110101000101001111011111110010",
8 => "011111011000111111100011101000011000111100101101110011011100010011110001110011001100101010010000111111101100000000100110101100110000110000000100000100010010100011100001110111011100001111010110110011011000101011010001100110000000010010111101001011000000010",
9 => "101111011011010000101111010111101110101000101111111010111101011100001100101010100010010000111111010001001000000100111111010011111011000110010000011001111100111000111111001011111011100101100010101111100001100000011110001011100001011000111010100111110010110",
10 => "101011011111011010111101010000111110000000101101100011011000000110000101010100110101001000011110001100000101100110100011001111011011111010001111111001001000110111001001101011010110111001111011001000101011010101011000100100011000000011010011000010000101101",
11 => "101110110001011000010011000000000100001010001010101101111111001011111000111010101001101110111000111111000111000000001010000111111100100000111000101101110010101100001110100111000100011010111011001110010101000010011101011100011001101011110011011100001000100",
12 => "110000110101000010001011000001011010010110000101001010010101000010000000010100011010101100101010010111000011000111010001010101011010010110000100010001011000111110000101110111000101001101100110001101110101010111100111100111001111011010111010101010010111101",
13 => "010000011011110101101100110100110110100000101001101000010000001101000100000101101101101010100001101010011001011111000100111001101000001000110101000001101011111000111000010010100011110001011111011110010000011111101110100011011101110101000001000100111000010",
14 => "100111001100010000010011100110001100000001111111010001010111000100110110000001110001111011101000110001111111101111110001111001101001100000001011100100111100101101100100101010011110110101010100101101110100001011010010110110100100000111110101000001110000101",
15 => "101111100100111011111111101111101110101110101001101001111111001010111000101100111110111101010101010011010100000000111100101010110001101101111111000000101111010110001101110010101000100111111001001000000100110110101000000011000110110111100101101011111011001",
16 => "000000100010101010101010111101000010001010001110011011110000000100000100111001100000001111001100010011110001100100111000111111101110110001110111000010111110001100101100110011011000000001010001001010000110001111100011110100011100011001001000100100101010011",
17 => "100001110010111011110111100001110101011111111111101100111000010001110100110001101000100100000001011101110011000011011000000100100110001110011100011010111000110110010110110100111101010001010011111110101010111010111111011100001110101010100100011100000010011",
18 => "111110101100111001100101111100110011001110000110001011000010010011010001011101110110110100011101100011101000011111110011011101010110110011011011001000100011010111110101101101101100000011010000001010011100010010001000000111000000001110101110001011000110110",
19 => "001111111101010000000101001100000011110110100000000000011011001101100100111001001111111111010110001111110100111100101010011101000001001100100000011000111101010011001001010001100110111101101010010100110001010001111110011110011101110000101010011100101101010",
20 => "100010000001101001101000111100101111010000010001010011101000011100111001100100111010101000010001110101111001101100000110000100101001111000000001001110111001110111000100000000110100100110100111001011011101111001111100000100100111101111100110001111110001011",
21 => "111010010111101100111111100110101000100011111100011110111000101000101100010001010001010000111001100010111111000100000010101011111011111001010110001000000101111101110000000101011100101111111101001011101111100111110010001110000000001000011010100000001110011",
22 => "000100010100000010100111101011111110011110000100000111100101011000011111110101100000001111011010101111001011000111101101111000110110011010100101010011101101010001001010001001110001111111101101011110110000111111000001111100100000001111100001110111010000011",
23 => "110000010111001111111100101000111011101000110000110111000110110000101011111111011000000000101111100101100110000001100100111011101111001110011101111000011000100111110111100011000011010100001011010000011010001111100101001100010000101111010110011000001011010",
24 => "111110000000011001011000111010000100111110010001101111011001000101001110000010100110001100110000010010111111111111110010101000111001101111010001000001111001010101001011001111100000110110000000101010011010001100101000000101101101011110111011100001000010100",
25 => "111101111111000100000010100110101000110101101001011111001010111000001010011100000101111010101000000111110010100110011010100010111001100100101001001111011111010100100100011010100001011011110110001010111111000010111000100110000100001011111000101101011010000",
26 => "100010100000001110011000110010010110011101110100110100100011111001011100000011101001011011101110110001001010010111110100100010001111000101010000001010010010000011010110111001110111100100100110011001000010110000011001110100100110111001011101001000101000010",
27 => "110001110000001011100101101111001100110101010010011100101100110100110001110010110111001010010011111110110110100011000001010010100011111111010110101010110011100111101110100101000101100110111101101110110100111010011011010001111111010101110111111000100001110",
28 => "001001010011000011010000101100001111001011100001000010100001101011111100100000010100110111110011001000100101010010000011110011011101111101010110001101000001111100101111011001001111110010000001101001011001001101001110010000010010100101100101011001101111111",
29 => "001011100011011100001101010011110010011001111010001100101110011111100010101000111010101010100100111101010111000011101000001101101010100100101011001001100000111001111001111100001010101111010011000110110100111111010001011110110010101100110011111011011110001",
30 => "011010011001110010000011000101100110101101011100101111100111010101000011000101001110100000000100111101000100010111011000101110000100010001110101010101011110110001011010100100111100010110010001010101010100101110010010001011111100001100011111001010100101110",
31 => "010101111111000010000101111001110111011110101001000011111001101110111001101011011101011100100100010010111100001001010011111111101000100100111111100011111001110000011101010111100010000101111101011000110100111010100111100001110001010100100000100101001010001",
32 => "110010100110010111111101000010000000001000000111100011010000111101010110111101000011001101000000010000010111001110010001001101101010011011100101110111100111011101010101100101101101000100101101001101011101100001111101110011001011111010001010000011110100001",
33 => "111010101100101110001010011111100100101000000100000001110110101011111100001001110101111100001001011000000001011000001111010011110110101110010111101001110110111011101010100110100111011110111000010011111001001110101000001110101011110011010001100010110110010",
34 => "011110111001110110101100101000010000001101110100001001000010000101001110000101000010000000011101011010000111101110000111100001000000111101101111001110110011011110110011101011001101010010000001010001101011001111111100111010011011110011111110011101001011000",
35 => "100101001010101001001101011111101011001000001000101100010010110010101001100110100000000000110011010100100101010000111111001111100101101011100000101011110100101001011101011100110110110110100100111111000100001111101011000000101101110010001010101011001010110",
36 => "001100011011000111101010000010001010001011110000100000100110010100111011000011111010010010100100111100001010111011001100110000100000000001100011010101001010100111100000001010111001101000100110000101001011001101100100001101000110000010110001001011111111101",
37 => "100001111101011110000010111011011011011000100101011101010111000101100100100100100101100110000110101101111010010000001000101011000000100111100010101100111110111000100111000110110100001111111001001101100100000000001100001010111010100001010101110100101101010",
38 => "100000011101010001011110101001001101000101000010001001011001000010110001100001100101000011111011010110010101001000110101000101100001010101001010011010110001100100110010100000101000100000111011000001110011011010000010000000100111011110001010000110110001011",
39 => "000101001011010000101000111110001110011111001011111011100011011100101011100100111111101000111001100101101001010011010111001011111100001110100011000100010001111100011000110100101010010000001011111110011100000010011011111110111011000100100010100000111110010",
40 => "111101100110011011101111011000100100000100101111000001010000000101001000101110111110000100001011000111010100111001001010101110101000101110110111101100010110110000011011001100000111001000001001011111110000100001011111000010101111110000000011100111011111001",
41 => "001010100100101000001100000111111101000011010001000011111000010100010010000000100001011111011111111101011101100010010101000101010010111110001001011010101011111011000000111100101110100010011001101101011011000000011000101110100101111100101110101000100000000",
42 => "010100010110101011001100001101010010001111010000110110010101110010101010011010010111000001001100010110110101111101100010001110001011101101101101100111011000000001110101001011011100100111100001110001000100110010000110011010110010110010111011111101001001100",
43 => "111100100111100110110101110000001101100110011001100110101111110111101000100111111011010110010001110011000101000000010001001110101111000011110001100010111000111111111001010010100000011110100010001010111001001100111000001100110010101100101010110011110010111",
44 => "000000000000010010100111011001001100101110100001111100110110010101010111010010010110010101000100000011001001101011000100111101100111010010110101010101011111001111010010010001011101110100010100001011010110010110001110110011010100001011010101010011110000001",
45 => "100110001000111100010100110111011110101010000111100100101011111101101110101000000000000010001011101010011001000101001011010100100001000000011100011111000011010100101101001000111001111101011011001110100101000010011111000010110101110000000100100111001001111",
46 => "110100010101010000110111000100100101110010000011111001111010010011101111100111010000000101101001000001000011111001010110001011111010101001100001110100011001100001100101110101101111001101100011111010100000110101111101001101100001000110100001010101011101100",
47 => "110011011110111000001111011001001101000111100110011100000100100010110101101101100000100010010100100000011001101000011100010011110101010001110110100110010111000111101000010101110010110110100010011000100001011111001001001000001010000000110101110010101110010",
48 => "001010110100010000000011010101110110100101100111101110100111000110000010000100011000110010010110001111011010001010000101001010000110100101100010000011011010010101100000010010010001101000110011001110101001111100001011111000110000000011100101110111000000001",
49 => "110000000000001111000011111110011111110110111110110000010100110101110110001111110100001110101101111000110010000010010011000111100000010001001001010100011010110101000110111101011011100110100011010011110110000000010100110101101010101000010000001111100010111",
50 => "110010111111001101111001010111100100001011010001010011110110110011011110110001101010010001011100000111110101011100110101100100010101001010001101001110100111001101011101001100111111111000000100001000010010101111010000101100001100100010011010010010101011001",
51 => "111010101010110000011011111000001001010011111011010111101100111100011011010011100001110011011100110011110101110011001001001000111011110011100000001100101001000000001001011000101100011000100110100100010001110101001010110001110001100100011100110001011110000",
52 => "000000011011101111101001001110100100110110010110010101111010001111011010111101110100111010000111100011011010111111101100000111011011000111101101101001010000011100001011010101101010000001000000011111010100100101100011010111100000100110101100010110001100000",
53 => "110010110001010010010100010101110110011011111101110001111111011011100101111011101100100110010100010101101101001011110100001111001100111011100010100010110111101000110110011000101000111011111001100011111001001110110010011001000110001000101101011011110001111",
54 => "000111011101000011100100101000010001001010100011101000000010100111100000000011000110111011010010001110000011101000110010100000000001100000001010111011011110000111000111111001010100001000100011101011011010000000101000011111010011100001001011111100101100101",
55 => "101000000000010011111100110001111100111001000100011000111000100100101100110000101011111000100011000011101011101011011011101100010011000111110111101111111111001100010101011100101101010110010001010111011101100010000000010110101011111101100010100101000101100",
56 => "110010001001101010111101000001000011100010000010100110000000010011000011010001001011010011101000110000101010111010101000010101111110101111001011011110001111001110101010000101110101001010111111011000100101001111100110111111000001101000000110001110011110000",
57 => "010010111001010010100010101000101001011110011100001011100111100001111100111101110010110001101101011010011001000111100010101001101111101001000100011100000111000000110000000100000100101010000100101101011100100110011010001100110110010101101111110001010010001",
58 => "101001000110101011011011000100110010011111111001100100101011010010000000011101100001101110000101111111101010100111100101000001000010001100010001101001100010101001000110111110100011110111000111111101000010111101010000010101000010100110001111100010101101100",
59 => "111111000011101000111111001101010011101100101010111000110001001011010000001000110010101010101101010010100100110110101000101110110111110010100000111101110000000110000110000110110110011111001111010101000001111111100111100101000010101001001001011101111101111",
60 => "010110101100111000101110111001111011011110111111011101000101101010010000010001010010011000110110010100111101010111101010010011000110110000111111001100010100110111100001110111001100101100010101110110001010001010010100010111111000000100001111111000000001001",
61 => "111111000101100100010010101000111001101011101010111110001100100101011011000101111000010011010011000001010001101100110001100011010110000011111111110101100100100010011001111111111101000001000110011011010010100111010110000100111000010001011000101100000001010",
62 => "110001010000111000100111110111111000010100101110111111001000110000001000100111001110011100110010111100010100001111011001101011101101110011101010011011000100111001000101000011101001010001111101010001101100011000110100001010110001110110010000001100101010100",
63 => "011100101011000001111000101001001111000011110100010001101000010110010100110111001000110001100011101000011111000010011011010110000001000111101100011010111101001110011010001111110101111001110111100010100110011110000010011111001010000110011010111000010010011",
64 => "001001001110111000111010101110010101000111110011110000110100111001100010101100101011010111001100010101011011101001101001000111110000101101010001001000101110110110110111110110010000010011101001011111001001000000110101100110000001110110010101111011001110101",
65 => "001010101101001001100000110111110111001010011010111111101101100110011101110010011010011100100110001111011110010000010001001011110010100001110110001110011011011101001010001000001010011011101100111110110101101010101011111001100101001001110101010111101000000",
66 => "101111111000110010101111101000101100000001111111011100011101000101111110100101110110110110110111001010100010111011000001100110011111010001000011010111111100010000111010000101010101010011111100011111100101010010100100111010001000010010001110011000001011101",
67 => "101111100010001011001001000001111000111111110100011011100010101011111011101000100000000111100110011010101111010001001011000001001110100100001110010000100001101001011111000001101010101010110111101010000101111011010101101101011000110101111011000111111011000",
68 => "111001111001110011001011110010110100001000110000000101001100011011011001011111000100110010000101011111111010100100100000110011010011101100111111001011000101101100100000100011000110101101000100001000010000000000001100011110011001010001110101001001100111101",
69 => "010001011101000011000100001011011110111001101110001001010110101010111001001110110111001101100000110001100010010001010111101110000101110100111001101110000000010101101001010011011001001011110110111010011010011100001000111101000101110001010011100010001011001",
70 => "111100110110010101000010100100000010000111011010101000001100100010011101110100100101110110110101101110000010111101111111011111000110000100101011010010110001011101101000100010001010000101000100101100010100100101010010010100011000101101011100101100010100010",
71 => "011100011101010000101011010111111011100111111101010110011011100000010110000100111011110111111010000110101110111001010111100010110000001000001111001011010011000010010011100011110101001001010110001100101111010000010111010111100011011000000011100110001011111",
72 => "000010111101010101001011001100001101010111010101000001000010111011010001111110010001110110011011000000000101110000001110111011101010110110000010111001101111101110001110010011111110011011000100111010110001010001000100011111111101010010000010110101100101100",
73 => "010010010111011011001011001111000010111100111100111011010011100110110100100110111010100100011110110011111000100110101001000101110110101010001100001111011000101010000100011001111111010111010000111010000001010101010110100000100010100011000111000010010001011",
74 => "101011010101001111111011110011000000011100111010100111101111101110010101001100101100001101010001111111001010010001110000001011110001100100110100000111000101101111000001110101011011001010110010011010101110000011011010100001101101001101110101010001110110101",
75 => "100110101011100100111011011001110001101001001011001100000011110111001101010110110010101011011110101011100000011011001101000100000101111010000110011010111001101000111111100111000110010010110010001110100110010011001000100010110100101001111010111110100101011",
76 => "011101101000001010010011110001010011011100001011100000101000011000000000001001111101100101101010010001010111111010101001010001111111000101010111111100101000000010000110010011001110010100000100101011000000110001100110110011100010100110000011111101111101111",
77 => "111101110100001010101101011010111000001110100110010000010111010111000101100101101011100100010100001001010101110101001101100000000000111110100111001011001101011001101100100011110101001100000100100001101000011100111011110011011100010110010101100000110011110",
78 => "100111000010111100110000010001111000111100110111001101111100001001111111110110011010100010010010010001100001110011000100000001011010001101110111111000000000110111111101010101001101010110111011000110001010111000011101100000101110000011100010011011010011100",
79 => "101010111101011001100001101011000110001001110010110011000101011110110100110111011110101100110010011101011001010100010110100100110000010000010101101000000111110010100010110110011101110010110011001001011000000110011110000010011010110000100010110010000111010",
80 => "110111101111000100011111001111100000000011111000010001101101100001000100000100001100001011100100000111111010010111101100001101101010101101001000010001110011010001100110011010000010100101001010010001111010101110000000011011001110011100111010000110111001001",
81 => "011001011110000000111111111101101111101011110011000110101101100010011110010100001100110011001110001111100101111011010000111000101100101000110001111111000111010000111110111110001110100110011000001011110111111011111101110101011100101011100010101010100011010",
82 => "000110001101111110100101100101101110100000110101101000010101110100110000010101110000110000100110000010010111111100110010100111011011111001101110100100111010011101110111100110011000100100010000000000111010110011111111110001100010110110111001000110001001111",
83 => "001111110111101100001100101011001010010100111010111101001111010111100011011110111110111101110100010100001001011011000011100011101101111110001010001111010110000000100100100011111100000101011100111011111010001001010011001100001110100111010001011010000000110",
84 => "001110011011001010111010101001100010110000110000011001110110111111001110110101000001101101010111110001111000100100111110111001110111010111110100011110011111100010000010101010010111101011000001100010010011100010111001011000110000010010101001011110000100011",
85 => "001101101010000100101111101111011011000000110011001011101101010111111110000010011000001011001111011001100011100011011110101101011001001100111001111011000011001011101011110110111001011001011101101100011101110110110001010101100001101110001001101001110011010",
86 => "100010000000000100110001101010100110001101110001011111101010111111110000000100000010100010001111010001101100111001110001001001000001111011110001000010001110011001110011110111010101001100110100010100011110010110110101001100001011111100010011001111100001100",
87 => "110010010110010001011010000001110111100101111000000010110111011100010011011101101101000000010110000110010100101011111011101111101010100000001011101100010110001000011110000101110011011011010100001111011000010010111111001011011101010001101001101001010110101",
88 => "101111111000000111111000110100011101001110110001100001111010111011111011100110011110011001110001101011111111111010100000010111000000000110001000111111100101010101010010000011101110001011000101011110101000110001010011000110001000100110010110101100111110011",
89 => "011001010011101101110011001010100100101010101100011111000010010110111010110011110110100011100011100010100101001110101101111011110100001010101000111100011100101011001001110111010101010011111101100010110100110101011011100011000100001100001011101110011000011",
90 => "001010011100001100100110110001111101100111010111100101001010111110111000100111010100010001111010010001111000101110011110100011011001100100100100001000001101100101011110101110001000011110101111110100001100010010000001110010000110110111000001110010101100110",
91 => "111010101010010011001111011000011100011010100110101000100100011000001101000111101001100110110001101101000100101011101110000011101100011001010001100100000011000000101010111101101101100110111100011001011100110111110110101000100111110111101011001101010101001",
92 => "100110010011110001011000101100100001100000011100100100111000110101100101001100010100001111110001010011110110110001100011101001110110110000101001011001101000110010001111000010001000110001000110000000110111010011011001000011001001000000001111100001000001001",
93 => "011000110010011111101100101011000001011000110110110001011000001001001110101100001110001111110011110111001101111011101111110000101010001000100111111010001010010111010011011011111000011000111000110101000101000100011101010101101111101010010100110101001011100",
94 => "011011100110101101010110011001101101101010001111100110111010101111010010011100001100001110100010110001101010001011000010001100101010101010000001000101001000001110010011110111011110111000110010001000101010001011100000110010001111100010110010101011010010101",
95 => "010001001001001010111000011101010110111001001001001111110110101010011010110000100011001100101100000011000111100111100101110011001000111110010100101111000011010110001100000110111110010111111111110101000100110101110100101100000111111000100011000110001100100",
96 => "011011000000110011001110011010011100010101001101101101000011110011111110001110110101010100011110111111010000010111000101110101100010010110011001111111111010011000111111000110001101001011110011000101011001011001110001000001100101001101111110001001101101101",
97 => "001011110100000011100110101101000100010111001010011010101101110110011011001000110011110000110100011100111000010110010001001001011101111001101100011110100110000100110111011011011100000001000100010001100011011001001100111110110011111011000111000001100111110",
98 => "010000010111110001010100000011101011011010100001010010110000101111101000010010101000000101010011001111100011000101011001010010111010000000100011010100001010100001101110001111011000111110100100001100110111001110011010000100111110000111001011110000110000010",
99 => "011011000000100001010110011011010001100011011101111111010111101110110100011001011101000100010111010011100011110110001101000011111011001001010001011100010011111000001101110001110011001001111111011000101111010011010110010011001000111001110001010001011001100",
100 => "001001101010011011001111011011001000100000001001110100011000101001001100010011110000101100100010001010110101111100000010001111101011100110001110000001110010001111000000100100110010100011101100111000000011101101010100011011001111000000100000111101110111111"
);


begin

CLOCK_PROGRESS : process
	begin
		Clock<='0';
		wait for clk_period/2;
		Clock<='1';
		wait for clk_period/2;
end process;

tester : process (Clock)
begin

	--test <= ROM_R(0);
	--check <= ROM_C(0);

	if (counter = 100) then
		counter <= 1;
		test <= ROM_R(counter);
		check <= ROM_C(counter);
	else
		counter <= counter + 1;
		test <= ROM_R(counter);
		check <= ROM_C(counter);
	end if;

end process;


checker : process (Clock,result)
begin
	if (result = check) then
		ok <= '1';
	else
		ok <= '0';
	end if;
end process;


dut : Decoder
	port map(
		clock  => Clock,
		input	=> test,
		output => result
	);

end architecture;