LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

entity test is
end entity;

architecture test_arch of test is

signal testvektor : std_logic_vector(3 downto 0);
signal umm : std_logic_vector(3 downto 0);

type ROM_type is array (0 to 254) of std_logic_vector(7 downto 0);
constant ROM_alpha : ROM_type := ( 0 => "00000001",
									1 => "00000010",
									2 => "00000100",
									3 => "00001000",
									4 => "00010000",
									5 => "00100000",
									6 => "01000000",
									7 => "10000000",
									8 => "00011101",
									9 => "00111010",
									10 => "01110100",
									11 => "11101000",
									12 => "11001101",
									13 => "10000111",
									14 => "00010011",
									15 => "00100110",
									16 => "01001100",
									17 => "10011000",
									18 => "00101101",
									19 => "01011010",
									20 => "10110100",
									21 => "01110101",
									22 => "11101010",
									23 => "11001001",
									24 => "10001111",
									25 => "00000011",
									26 => "00000110",
									27 => "00001100",
									28 => "00011000",
									29 => "00110000",
									30 => "01100000",
									31 => "11000000",
									32 => "10011101",
									33 => "00100111",
									34 => "01001110",
									35 => "10011100",
									36 => "00100101",
									37 => "01001010",
									38 => "10010100",
									39 => "00110101",
									40 => "01101010",
									41 => "11010100",
									42 => "10110101",
									43 => "01110111",
									44 => "11101110",
									45 => "11000001",
									46 => "10011111",
									47 => "00100011",
									48 => "01000110",
									49 => "10001100",
									50 => "00000101",
									51 => "00001010",
									52 => "00010100",
									53 => "00101000",
									54 => "01010000",
									55 => "10100000",
									56 => "01011101",
									57 => "10111010",
									58 => "01101001",
									59 => "11010010",
									60 => "10111001",
									61 => "01101111",
									62 => "11011110",
									63 => "10100001",
									64 => "01011111",
									65 => "10111110",
									66 => "01100001",
									67 => "11000010",
									68 => "10011001",
									69 => "00101111",
									70 => "01011110",
									71 => "10111100",
									72 => "01100101",
									73 => "11001010",
									74 => "10001001",
									75 => "00001111",
									76 => "00011110",
									77 => "00111100",
									78 => "01111000",
									79 => "11110000",
									80 => "11111101",
									81 => "11100111",
									82 => "11010011",
									83 => "10111011",
									84 => "01101011",
									85 => "11010110",
									86 => "10110001",
									87 => "01111111",
									88 => "11111110",
									89 => "11100001",
									90 => "11011111",
									91 => "10100011",
									92 => "01011011",
									93 => "10110110",
									94 => "01110001",
									95 => "11100010",
									96 => "11011001",
									97 => "10101111",
									98 => "01000011",
									99 => "10000110",
									100 => "00010001",
									101 => "00100010",
									102 => "01000100",
									103 => "10001000",
									104 => "00001101",
									105 => "00011010",
									106 => "00110100",
									107 => "01101000",
									108 => "11010000",
									109 => "10111101",
									110 => "01100111",
									111 => "11001110",
									112 => "10000001",
									113 => "00011111",
									114 => "00111110",
									115 => "01111100",
									116 => "11111000",
									117 => "11101101",
									118 => "11000111",
									119 => "10010011",
									120 => "00111011",
									121 => "01110110",
									122 => "11101100",
									123 => "11000101",
									124 => "10010111",
									125 => "00110011",
									126 => "01100110",
									127 => "11001100",
									128 => "10000101",
									129 => "00010111",
									130 => "00101110",
									131 => "01011100",
									132 => "10111000",
									133 => "01101101",
									134 => "11011010",
									135 => "10101001",
									136 => "01001111",
									137 => "10011110",
									138 => "00100001",
									139 => "01000010",
									140 => "10000100",
									141 => "00010101",
									142 => "00101010",
									143 => "01010100",
									144 => "10101000",
									145 => "01001101",
									146 => "10011010",
									147 => "00101001",
									148 => "01010010",
									149 => "10100100",
									150 => "01010101",
									151 => "10101010",
									152 => "01001001",
									153 => "10010010",
									154 => "00111001",
									155 => "01110010",
									156 => "11100100",
									157 => "11010101",
									158 => "10110111",
									159 => "01110011",
									160 => "11100110",
									161 => "11010001",
									162 => "10111111",
									163 => "01100011",
									164 => "11000110",
									165 => "10010001",
									166 => "00111111",
									167 => "01111110",
									168 => "11111100",
									169 => "11100101",
									170 => "11010111",
									171 => "10110011",
									172 => "01111011",
									173 => "11110110",
									174 => "11110001",
									175 => "11111111",
									176 => "11100011",
									177 => "11011011",
									178 => "10101011",
									179 => "01001011",
									180 => "10010110",
									181 => "00110001",
									182 => "01100010",
									183 => "11000100",
									184 => "10010101",
									185 => "00110111",
									186 => "01101110",
									187 => "11011100",
									188 => "10100101",
									189 => "01010111",
									190 => "10101110",
									191 => "01000001",
									192 => "10000010",
									193 => "00011001",
									194 => "00110010",
									195 => "01100100",
									196 => "11001000",
									197 => "10001101",
									198 => "00000111",
									199 => "00001110",
									200 => "00011100",
									201 => "00111000",
									202 => "01110000",
									203 => "11100000",
									204 => "11011101",
									205 => "10100111",
									206 => "01010011",
									207 => "10100110",
									208 => "01010001",
									209 => "10100010",
									210 => "01011001",
									211 => "10110010",
									212 => "01111001",
									213 => "11110010",
									214 => "11111001",
									215 => "11101111",
									216 => "11000011",
									217 => "10011011",
									218 => "00101011",
									219 => "01010110",
									220 => "10101100",
									221 => "01000101",
									222 => "10001010",
									223 => "00001001",
									224 => "00010010",
									225 => "00100100",
									226 => "01001000",
									227 => "10010000",
									228 => "00111101",
									229 => "01111010",
									230 => "11110100",
									231 => "11110101",
									232 => "11110111",
									233 => "11110011",
									234 => "11111011",
									235 => "11101011",
									236 => "11001011",
									237 => "10001011",
									238 => "00001011",
									239 => "00010110",
									240 => "00101100",
									241 => "01011000",
									242 => "10110000",
									243 => "01111101",
									244 => "11111010",
									245 => "11101001",
									246 => "11001111",
									247 => "10000011",
									248 => "00011011",
									249 => "00110110",
									250 => "01101100",
									251 => "11011000",
									252 => "10101101",
									253 => "01000111",
									254 => "10001110");
									
									
									
type ROM_type2 is array (0 to 254) of integer;
constant ROM_alphaInv : ROM_type2 := ( 0 => 0,
1 => 1,
2 => 25,
3 => 2,
4 => 50,
5 => 26,
6 => 198,
7 => 3,
8 => 223,
9 => 51,
10 => 238,
11 => 27,
12 => 104,
13 => 199,
14 => 75,
15 => 4,
16 => 100,
17 => 224,
18 => 14,
19 => 52,
20 => 141,
21 => 239,
22 => 129,
23 => 28,
24 => 193,
25 => 105,
26 => 248,
27 => 200,
28 => 8,
29 => 76,
30 => 113,
31 => 5,
32 => 138,
33 => 101,
34 => 47,
35 => 225,
36 => 36,
37 => 15,
38 => 33,
39 => 53,
40 => 147,
41 => 142,
42 => 218,
43 => 240,
44 => 18,
45 => 130,
46 => 69,
47 => 29,
48 => 181,
49 => 194,
50 => 125,
51 => 106,
52 => 39,
53 => 249,
54 => 185,
55 => 201,
56 => 154,
57 => 9,
58 => 120,
59 => 77,
60 => 228,
61 => 114,
62 => 166,
63 => 6,
64 => 191,
65 => 139,
66 => 98,
67 => 102,
68 => 221,
69 => 48,
70 => 253,
71 => 226,
72 => 152,
73 => 37,
74 => 179,
75 => 16,
76 => 145,
77 => 34,
78 => 136,
79 => 54,
80 => 208,
81 => 148,
82 => 206,
83 => 143,
84 => 150,
85 => 219,
86 => 189,
87 => 241,
88 => 210,
89 => 19,
90 => 92,
91 => 131,
92 => 56,
93 => 70,
94 => 64,
95 => 30,
96 => 66,
97 => 182,
98 => 163,
99 => 195,
100 => 72,
101 => 126,
102 => 110,
103 => 107,
104 => 58,
105 => 40,
106 => 84,
107 => 250,
108 => 133,
109 => 186,
110 => 61,
111 => 202,
112 => 94,
113 => 155,
114 => 159,
115 => 10,
116 => 21,
117 => 121,
118 => 43,
119 => 78,
120 => 212,
121 => 229,
122 => 172,
123 => 115,
124 => 243,
125 => 167,
126 => 87,
127 => 7,
128 => 112,
129 => 192,
130 => 247,
131 => 140,
132 => 128,
133 => 99,
134 => 13,
135 => 103,
136 => 74,
137 => 222,
138 => 237,
139 => 49,
140 => 197,
141 => 254,
142 => 24,
143 => 227,
144 => 165,
145 => 153,
146 => 119,
147 => 38,
148 => 184,
149 => 180,
150 => 124,
151 => 17,
152 => 68,
153 => 146,
154 => 217,
155 => 35,
156 => 32,
157 => 137,
158 => 46,
159 => 55,
160 => 63,
161 => 209,
162 => 91,
163 => 149,
164 => 188,
165 => 207,
166 => 205,
167 => 144,
168 => 135,
169 => 151,
170 => 178,
171 => 220,
172 => 252,
173 => 190,
174 => 97,
175 => 242,
176 => 86,
177 => 211,
178 => 171,
179 => 20,
180 => 42,
181 => 93,
182 => 158,
183 => 132,
184 => 60,
185 => 57,
186 => 83,
187 => 71,
188 => 109,
189 => 65,
190 => 162,
191 => 31,
192 => 45,
193 => 67,
194 => 216,
195 => 183,
196 => 123,
197 => 164,
198 => 118,
199 => 196,
200 => 23,
201 => 73,
202 => 236,
203 => 127,
204 => 12,
205 => 111,
206 => 246,
207 => 108,
208 => 161,
209 => 59,
210 => 82,
211 => 41,
212 => 157,
213 => 85,
214 => 170,
215 => 251,
216 => 96,
217 => 134,
218 => 177,
219 => 187,
220 => 204,
221 => 62,
222 => 90,
223 => 203,
224 => 89,
225 => 95,
226 => 176,
227 => 156,
228 => 169,
229 => 160,
230 => 81,
231 => 11,
232 => 245,
233 => 22,
234 => 235,
235 => 122,
236 => 117,
237 => 44,
238 => 215,
239 => 79,
240 => 174,
241 => 213,
242 => 233,
243 => 230,
244 => 231,
245 => 173,
246 => 232,
247 => 116,
248 => 214,
249 => 244,
250 => 234,
251 => 168,
252 => 80,
253 => 88,
254 => 175
);

begin
	
umm <= "0011";
	
testvektor(0) <= '0' xor umm(0);
testvektor(1) <= '1' xor umm(1);
testvektor(2) <= '0' xor umm(2);
testvektor(3) <= '1' xor umm(3);



end architecture;

