library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.std_logic_unsigned.all;
--=======================================================
--  Entity decleration
--=======================================================

--DE10_LITE_Empty_Top: 
--
-------------- CLOCK ----------
--input 		          		ADC_CLK_10,
--input 		          		MAX10_CLK1_50,
--input 		          		MAX10_CLK2_50,
--
-------------- SDRAM ----------
--output		    [12:0]		DRAM_ADDR,
--output		     [1:0]		DRAM_BA,
--output		          		DRAM_CAS_N,
--output		          		DRAM_CKE,
--output		          		DRAM_CLK,
--output		          		DRAM_CS_N,
--inout 		    [15:0]		DRAM_DQ,
--output		          		DRAM_LDQM,
--output		          		DRAM_RAS_N,
--output		          		DRAM_UDQM,
--output		          		DRAM_WE_N,
--
-------------- SEG7 ----------
--output		     [7:0]		HEX0,
--output		     [7:0]		HEX1,
--output		     [7:0]		HEX2,
--output		     [7:0]		HEX3,
--output		     [7:0]		HEX4,
--output		     [7:0]		HEX5,
--
-------------- KEY ----------
--input 		     [1:0]		KEY,
--
-------------- LED ----------
--output		     [9:0]		LEDR,
--
-------------- SW ----------
--input 		     [9:0]		SW,
--
-------------- VGA ----------
--output		     [3:0]		VGA_B,
--output		     [3:0]		VGA_G,
--output		          		VGA_HS,
--output		     [3:0]		VGA_R,
--output		          		VGA_VS,
--
-------------- Accelerometer ----------
--output		          		GSENSOR_CS_N,
--input 		     [2:1]		GSENSOR_INT,
--output		          		GSENSOR_SCLK,
--inout 		          		GSENSOR_SDI,
--inout 		          		GSENSOR_SDO,
--
-------------- Arduino ----------
--inout 		    [15:0]		ARDUINO_IO,
--inout 		          		ARDUINO_RESET_N,
--
-------------- GPIO, GPIO connect to GPIO Default ----------

entity Encoder_Top is
  port (
		KEY        : in std_logic_vector(0 downto 0);
		SW         : in std_logic_vector(0 downto 0);
		ADC_CLK_10 : in std_logic;
		LEDR       : out std_logic_vector(7 downto 0)
  );
end entity;

--=======================================================
-- Architecture declaration
--=======================================================

architecture HWTB_arch of Encoder_Top is

	component product_encoder
		port (
			clk : std_logic;
			rst : std_logic;
			X   : in  std_logic_vector(238 downto 0);
			C   : out std_logic_vector(255 downto 0)
		);
	end component;
	
	type X_type is array (0 to 238) of std_logic_vector(238 downto 0);
	type C_type is array (0 to 255) of std_logic_vector(255 downto 0);
	
	constant X_data : X_type := (
	000 => "11000100101010111111010011111001001011010111101011010111010111011111010011001000011111100100011100010010100001000100111101100111111101010101110100111100110010101001101101101001101110011110100001001100001001001000111011110110110101001001111",
001 => "10101001001111001101011101111111110011001010001100011100111110111010110110010100100001011010001101110110011010001110011001111011111100110111101100011101110001000110000111010000011100101010111001011001110010110011000011111101010110000100111",
002 => "00011110101101111011000001011001010010001001111010010001101100011101000011000011111011001010100101110001101000111000101010110100000000001101010111110100011010010000001111110110100001011010101011011111101110111101100011101000110110011110110",
003 => "10011110000100100101110001111111110111010111101100111110100000001011000001010111100111011111011111110000001101101000000000111000101100010110011101001111001011001000001000010011001010000000011011101110110101000010001100100110111000000000111",
004 => "10011111100101100111000100111011001110001000001011110010000000101111101001100000110001001000110001001011100100000110101000100111011010110000100001011001000011001101001111100011010001001001000111010110010110101011010001010111110011011101111",
005 => "10010010110110100111110110000010100100101001101111001000101000111100110110100000111001000001101011000100100001100011111000101011011001101011100100000011111011110001001110111011110000110001010100001001010000001111010100001111000110000100110",
006 => "01011010101011010001101011010110100100101100001010111100100110111001101001011001001001101011010111000011100100000000001011100001110011110111011000110111011000110011100100001010101111110001000001000111000000000000010111010010101111101001101",
007 => "00000011101011000110010011011110001011100001101000010100011101010010101100111111011001111010000010000111000010000010101010101001011101111010100110010110011011100010101110001001001100110101011111111111011111100010101000010100010010111000000",
008 => "10001111110110000000111011000000100111111001100011010110110001110010110011011010110111101001111110100100010010110100100000001011011111010111010000100011110011110110110110001001100101111011011001001011110101001110101000101111011100010101010",
009 => "10001010101101001101000101100001100010111001011000110100111100011111001011101010111100010010011110010000111111010001111110010001110100011000111000001110100000101111000010110100111101100000001011110010000101010001000101011000000010010000100",
010 => "00100101111110000000110110000110011000001010000110111000100010011001001111011100000000101110100100101101110111110100001110111011110000011111100101110001000001001101000010001111100110000011010000010100111111111001001001111110100100101001110",
011 => "00011011001101101110111000110001010001110111001010111100001010100011001010001001011011101000011110001111001011010100111110110101010110010000110011001111100011101111011110001010001011100010000111101100111011101110001000101110110110001100101",
012 => "10101101011111010000100011001010001010100001110110010001110111010001000001010101111010111100010000110011000110001101001110100110001111111001000010001001110010110100011000000100100110001101010100010000010110010110011111011111001101111111000",
013 => "00110000010100111111010011000011111100100101100010110010010000101111110010100000101111111001111100000000110000001011111000111111110001100100111000001110101010000100100110000001011111100011010001011000100111000010110111111011101001111010011",
014 => "00000001010010010111010101011100110010010101000111010110001011011100011101011000111100101010101010100011100100100001010110010100110010011011001110010101000111001111100100000100000100111110011101001000001101101001010000110111100011010010110",
015 => "10111101010000110100011110010110101011101001001101011000000000110111010010011101010010111001001010100100110010001011101101001010111011110111101100100100011001001100000001101001100000010101110001111110101111000101010111001010110101001111001",
016 => "01000110000111111111001010001111111100111110001010001011111101010001000100010011100011011111111010010110101001100001100000110011011110100001000011000100000011111011010010011100110111001110000000010101000110100011100000011001111001001011001",
017 => "11011010000111000001000111100101111101110001001110111101110111100001001100100000001101110000010111101011011010001101101110110000000100111000101101011000001100110000110010111001001011001000011101111100110111001100000000001100110010100110001",
018 => "00110101000111000101111011101111010101001010000001110001110010001011010101110100100101111011000010101101111100000101011010111111100101110101010101101111100010110100110101011100011101011101100000110101110010101110100001011001001111010010100",
019 => "00001110011000100010111000000000110010010010100110101100011100101111110010110011100101101010000101010110001110011111110000010110000100000001100111111101011101110000000010001001111001101101011011111111010111111010111101100000011100100000110",
020 => "01010001110100110001000001001010101100101111001010101010001011010100010101001100010010000000011010000001010110111000010011111010100101110001100001000111000000100010010011111111011101101100100101010011100110000010110011110011000101000011010",
021 => "11000010000100110100011000111110000011000010111110011011000111110000010000011100111101011011000111111000111011100101111111000110100001010111101000111100100000010101011101010000011111111010001110110001001100010000111101101110010000101110011",
022 => "10000001100011111011011000101000110101010111011110011001000010110110101111110110101110001111100000110110111010100001000101101101111001101011101001110011011100001011100111111010110110010111110110101101001111111101110011111000110101001110100",
023 => "00001110001011101011100100000101010001011100101001100001100011001011101001111010011100000101101110010001101110001000000101000100111000100010111010111000000111010000001101110000010001000110001110011001101001000111110001110011110001000101110",
024 => "11110101100110011111110010011001110100001100000110011100010110100100001110110011100010001001010011100111110111011011001100010110001101111101110100000101101100100000111001011001100010010110110011010010000111000101001001111110111110100101110",
025 => "11001000101100010101101111110001010000010010100011100101111010010011001001011100001100110100001110001100011010010010001111101001110111110001011100000101011001000101001001111111111101101111001001011011100110001100010110111011110100000011010",
026 => "10001111011110010010010010111010111101111111001101110011001011001000001001001110000111101100011111101000000010000000110110011011000110010010000001011100001011001010101000110111010101111111000010011101111011011111101101100010011001100010110",
027 => "00101011001010111000110001111101010111110110100100100010111110100111000110010011100100011011101101111111000000110011001011101000011110111111011010101110111111001001000011111011100111101001111110101100011111010011011010101001100010101110101",
028 => "11001100011001110110001001100110101111110110011111001111001100001011000100000000000111001111001011100110111110100110101000011101111001110101011111010010010001111110111110111100000110001110101001100011100100100111111111111000111011101101100",
029 => "11101111101000110010010000010111100101011111001010000111100101100001101010111101101010110011101110000110011100010100100100100110001011100101001001101100111010010110110000000101110001000110011000010100000111110010000111010101000011000111100",
030 => "00101100100101001011110000010111000101111011000100011100111100110000101000000010000000011100011001011010101100010000100010001010100000010110100110110011111000010001001000110001001011000100001110110000101000011000011111110100000000101110100",
031 => "10110110111110001000001010001111101100000001100010011100100010111001110111110100101111011101110110100011011110110110101110110001000011111011001111011100000000100010000010011011011110011110100110010010111011000101110011011001100011100011111",
032 => "11100101111100100011010001001100101111000111010100010011110100001111010101010101111110010100001000000101000001100010110011100100010110000000110111010100011010000011101100000001101001011111000111011110111100000000101101110011011100101001010",
033 => "10000010010000000111101010100011000010011010111010010000110001000010100110001000100110000100010000000011100111010000100110011000001111010001100001000110001110110010010111100110111110101000100111001100000011011111110010100010111011001101000",
034 => "11110000101111011111010001101001101011101001101100100010001111111010110110110010111110011011110111000101001110011100110100010100011001001010101000100100100100111110111101000101011001011110011011101111010000001101011000101101001001101111001",
035 => "11100011111001101101001101001001000100011100101100011010100010111000101011110000000111100010011010000001110001011011110100110100100010110111101011000101110110011101000000011010001101011101100110011111011010000100101111010111110001110101011",
036 => "01101000011100111101111010110011101101000010011001010110011100110110001110011001100111111110001000101011101001100110001110100100010101111000101011011000101011111101100010001100001011000100011110111000010110100100100001010011010100000011010",
037 => "01010110101000110000110001101010001010000010010111101101010001111101100001000100010111101101011001101001011000111101111111111010011111110011010110110010100101010100111101111010010110010110100010000000101011100100011100111000110111110011000",
038 => "00000111100011011100100000100101111100111101111110010111011001000100010101010110011001110111010110000001010100101001001011111101011100011000100111010010011011111101100011010100111001111000011111000010111000100011110001001011010110010110101",
039 => "01111001000111000011110100110101100011111001001001000111111110101010100111101011101001100110101110101111011011110100001011010000111000010100001110001111110100000000010101101100010100111001010010100000001010111000010111010111011000000100111",
040 => "10001110000010111110000000010100001001110010100010010110101011001110011101001110100110011011101010111111001000111001101110010111101101100000010010010001000110111100001101101001001001101111011010010101101011100010000110000000111100000010110",
041 => "01101001001011111010010111010100100011100110101011110110001010001010110001001001001111100111111101000011001001000001010110101001001001111101001011101100011011011000101111100101111100101111110000011110010111011000001001010010111101010000100",
042 => "11110011010110101001100001011010110011011101010110111110111111001110011000110100110000010001001111101011101111100100000011010101110100011010011110101010101100111101101100010101010000100111110000111001101010011010000001011111000111010111111",
043 => "01110001001100010000000000101100111000101000010001010010011101101101000110000100010011010100101111011001010100101001010011001101111000101011000100101011010100001010010000101111101001001100001110101111111010110001001111111011011011010010111",
044 => "00101111011011000100011110101011011111100011011001101000000011111100111100100000100000100101111001110011100101001111111000011001000001100100101111011110001111110011110011111110101101100010101010100101001111001111001111110100011100110011010",
045 => "11011100111011100100110110101000101111100101001000001110110110111111011111101011010100110010111100001010100011010100010111011010001000111111100111001111000001010111000110110010111110000110110000111110100000100000110100000010001010001000000",
046 => "11000110010011101000101010100110100110101010101010110010001101000010101001111011000111110010110101011110010011110011101001010011110111111111111111000110100000101101001100001110100000111010001011010101110100101110110001010111000010110011011",
047 => "11011010111010101000000011000010100011010011001011010010011111111111110011000001110100000011110100010001011111010111110100001101011001111000011010010100111111000011000110101001111101001111111011111110101011011000011011010011110011010000010",
048 => "01001000011000011111011111100100100001111010010110110100010010101110000101000100010011000010100111000001000111001001011111101001100111110111101110011111000001001000101011110100110110001011110011000010111100001011011010001111101101000000110",
049 => "11000111010001001111011110011010010010011000100111001000111001011010101000011110111101010011100101011010100010111011100000110001101111001101010100010011110010111111001110010111010010010111001010001110001000111001101110000101010101010101111",
050 => "10110101110011011100111110101101100100011001011111111000101000100100100110010011101100100011111101011001000011111010010110001101011101101111111001101110110010100100100010100111001010100011001110111101000110101000101100001000111010010111010",
051 => "00010110011000110010110000001111111000101001001100111101010100100110101011111110010101110010110010100001111111110001000000110111100101010100101101000110010101011011100111001011111000000001011111110100111011111100100111111001000110010111111",
052 => "11011001001000001110111001010000010111100010000101110001011011000010100010110110010111101111110111111011010111111111010101011011101100010011000000000011110111010001111010001000001011101110101101100011101100011110011010010000100010111101010",
053 => "10010100111010010001001011000011000000001101001001110001111000001111100010100111100111011010000011000000111111110111111110101111011101101111001010110101001001001011101101100010101111101110100111011101111101100010110101001001001110010010010",
054 => "10111001011011010101101101110001011100100101011100011001111001100110011000001101001011101100010101000100011001000110011001100110001000001011000010111000011000001111101010100100110101000010111100010010000010110000110110010101001001000001111",
055 => "10111111000101010011100100111111011011110011110100100010110011011011010011101111100100011011000011011101101110101111011000011010011010100111001110110010001111010110001010100111110001010111001001010011101010110001100111000011000000101011010",
056 => "00100011101101111010100101000111010100100111110110000011111101011111010100111010011010011011000110100001101010101111100000111011101100010001101000110001110011111010000110111110010100100101001111011101010000000100101100001101010101001000110",
057 => "10001111110010001010100111101010101110111011110001111111101001110111010001011010010011001100011001101010111010010100011101011010110010010000010110000011100001001100010011100111100110010010001011011011111011011110110011011000111011110101111",
058 => "00110110111111001101101000001000111100000110111001011111101011010010110010001000110010110111010100100110011000100000000111001000110010111011011111101001000001001110010101010011100010011111110011010100000001110111111110110100110110100110101",
059 => "11011001100011111010010110110101111011101100111000100101111010010011011010010111111111110100010111100011100111010100001110000011111101110000000010000101011100011001101111000001101000011010110110001100010000011110010100001110111011110000011",
060 => "00101110111001001011001111111111000100101011011001011000011011010000001011100000101010100001011011111000110010110001000110100100011011100100010000000000011100000111111100110100101110011001111010001101111011110000101110010011110101000010001",
061 => "00001010110010101100001101001001101001001101000101000010010101001011110010011000111011001010101000101011000111110100001001001111001111111011011101011100110100101110010101010100011010010011101101011111110100100110100001101001011101010011000",
062 => "00000001001100011111110000010001101110000010001000010101001111011011111110101000001111010100000010101111011010100011000010111001011100001000110000011100011000011010011111101101010011010000100010000111100100101001011000101011010001111000100",
063 => "00100001101110100001000110000101000010010111001011011101111111111111111000111010100000010110110011000101001000001101111110011000010100000110001000010010000111001001110101010010011011011001100110001110000110100011110010010001111011110001010",
064 => "00100010100111001101111000011100011010101100110111001111001110100000001001100011001110111011110011110011100100101001010000011100111000111011111111011001111000101011000111110000010001100011010010111010010111100001100110000011110100001100111",
065 => "01101010010000011001010010111111111110010010111111001101011000001100010100010001111010101010000000001110001111101110111100101101010010101001110010110101110111010010110110111010011111101101000111100100101100011100010000001010010101011010101",
066 => "10001101111100100011111011111110010100110100110101001000011110101110110000110001000000000100001110101001110001100100110100111101000011101111001000000010111100000101110111001001010010110011011110100000001100111111100001001101100010011101011",
067 => "10111010110011000000101000101001011111101000010101110011000011101011001111110010001100101111010100001100110010000111000110110011010111010001110100110101001001010010010100111111001110000001010101101111111001001001101101111011101011010100110",
068 => "00101001101111000010011110000111001011100010110001101101001001101100111101011110000101011001001111101001110101010010111111001000110001101100101101101110000100111011100100100000011001000111010100001110010010111000101101101001111010001001110",
069 => "00010010111101110001111010011000111111100101101100110101100110100000111001000100010001101101000000110011010110111001111010110110001111000011101001111100001110000010111111011100110010100110100000000101010000011100011110011101001010011111101",
070 => "10110011000110000101101011011100010101011010000010111111010111101011011111101101001101110001100011000011110000111010000000101011000101000100111101001111101011011001010100011101011001111010010110010100111011010011011100111111110000101110110",
071 => "11101001010100001000110001100010010010000110001011011000010110101000101101101100000010100111111111111000010110100011000000000000100010011011000100000100000111101001011101110001010111010010100000110010101101010010011100000110010010010110110",
072 => "00111101001101110000010001100101010011111111001101010011010000111100011111011000101101111011111000001010110011011011111101101001100100111001001000111100101101101101111001001111001011111001010110010111010001000011010111101011111111000010111",
073 => "10010110011101111110011100000010000101011100001110111110111010000111100110001011101100001101101000001110100101000101101000100001001010010100000100110101110011101000000101010010110111110001010100000111100011110010010111011111010010001110101",
074 => "00001101011110010111100110001001000000001001111101101100110001110100101011111000110010000110110110001001001000100100100011001110100110011000000011110000100000101001010100101001101100010101011100100001010101000011011100110111100001010100011",
075 => "10001100101100100010101101011101010000110011010011100111011000010110101111010101010000101100010110100000100101110100101000000110011110100100111010000011101101001101001011110111100011001000100100011010110110111010110110000100110100111100011",
076 => "11111000011100101010101011011111100001010000010010000010010011110101111101101100011101010111100011100110011110010110100101111010100010011100010011101011100110000001000001010100010110110010000110011000100101001111011001110011000001000100110",
077 => "00010101001011000111101011011101001010010100010001111011110100100101011111010000010110000101000001001010001000101101000100111101100111000100001111011111011110111111000111010010000000100100010100101001001011011010001011011011110001000011100",
078 => "10101011100000011100101010010100000010011011111010110001000111110101000101110110010100001111111010111100000001001101011000010100110010111110000111111110111110101111110101000100111110111100101101010110111101011111100101010000101000001111100",
079 => "10110101111101001110101001001000010011101111000100110000100001111000010111010001111010010001100000111001000011101100100111110100101010111010100011111110110100010101011110000110000010010110100101111001000001001011101111110001101101110001111",
080 => "11001110111010001110001010011101110100000000100000100110001001111011010001011001101110000000101111100110000100100100010011010010110100111101101111100000100100011011010110110001001000001010000000011110111101101010001011001000110001100010011",
081 => "01000111011100111000010111000100000001111010001111100101000000100000101001000110101011010101001000011010000111100011101101010010111111001101001001000010111000011011100101111000010010011100010000100100000111001100000010011001101011011100011",
082 => "01111101100111010011101010001101110101111110010100000101100110011100110101100110001000100001001101011110111101111000110110100010111111100101101011100000011010010101010010010001001110110100101111100010011111101110001001000001011111011111101",
083 => "10110101110111011011000110011010011011001010111101101001110001101000011000001110111001000001111010001010110001101001001000010101000100010110001101111001000100001000101101110101010110001001111010101010110111001100000011011001101011010001100",
084 => "10110100111001101111011101111110110100111110000000100101100101001011010010110101100000001100011111111111010110110000111111000011000001011000101101100100001010010101101011110011011000101110110010101100100101001111010011000101100111101001010",
085 => "11010111010001011110111001111101010100100111111110101010111111111010011100011011110111111000011101111101001101010111001100001001011101100111110110011010101111000110110001010101111101000101100101101001001010111001000100010001111011110000111",
086 => "11110110001101010010101000110000001111010110110010000011011001001100100110011101011000000101100100000100100110011100111111101000010000111110011101010001110010111100111010010011111100010000110100010011011101110111011111011101010011010011100",
087 => "01100011010110010001101100110100011000001001011011010000111100111110001000101100011110000000110011100011101101011010011100111000011000000011110111110011101100000010000011011000011011000101100011011011000101101001110100110011111000001011010",
088 => "11111011011001000100010010110110001011101110010100100110010110001110001010110010011000010010101100101111100110011011101011000100000001011111001011111001001010001010110100010011000011100001011011111010011101011011001110100001101101100100001",
089 => "10111101000000011110100100001101000100111101101111001001000000100111001010010000000001000110110010111101010111100100011100100110010101110000010001011101011001100001010101101000000001000111100110011010010001001011100101000001010011011001011",
090 => "10011111011010100001011000110001010100101001100100111111100101101101111110100111011100011010100010110101000100101101001100001101101001001000110111110010101101111000001011100101010000110101101011000001110001100001100011011000011001111100111",
091 => "01010100111110101011100000111101100010110010110000101001101101000100010010111000000100111000110101101100110110010000100010110100010011111100101010010111010001111100000110011100111001010111000101000100010111010010110110111110111001101100110",
092 => "00101001100101010001001011110100111000000000100101001001100100011000110101101111010100111011001110100101110000010011111111110010000001101010011001111101010010100000100111001110001000010010011011010000010101100001100010010001000011011110001",
093 => "01111101010101111111101010011110000010011111011011110011100010001101110010001000010011110111110010101011101000100111110110010101001110011011111110000010111010000011010111001010001111000011101101011101001010111110101010010001101001110001101",
094 => "10011000001001110100101101011111100001010010100111110101100101110001100100111111110010101101000101100010110010010001100011111000101101100100010100100101010101000110010011100010101000101001110000111000010111001111001100100011011110001101011",
095 => "10000011101111000000000000001100000010110110101011101011101001000001111001101101100101010011011011010000000101000111101000111011010101100100000011010010001001001001111000111101110101010011001010010010100111101011101111001111011000101011001",
096 => "01000110101000010010001001010110100110000111100111100111101001111110111001101111000011001111011111110000001101011100011100001001111111101110111110010100011000001010010001010000110111100001000100101001111000100110111011100100110010011101110",
097 => "10110011101010110011010010010010100000101000111100101101001111011000100011001000000110000000101111100011100110001101111110110111111010110110100110011101011110100100110101101100011110000101101001100101000000000111111010000011000001101111110",
098 => "11101100000101100001101010111000111000010011110111101010001011110111100100011010101001011001100100010001000110101000101111110001000100110001100011010101000001011110100010101111011000010000100110100010110101000110011101011001111100011111010",
099 => "11100000010101010110001011011011110111111110111111000010101001110110010010110000010010101011100000100110011111101001111001011010100100011111111111101000110000010100100100100101001001111111111011100011100101001100111011011100011000101010101",
100 => "10101110101001000010010100010110011011010111100010011000001011001110010000011111110100101001000010101110110000010100001101101000001111110001010000101001101101010101001101100011101101001011101100100001000110111010011110001101100101100011100",
101 => "00011101101001001110110000111011010001000000011110001111010001101001100010101010110000011110110101010001110000011001100000110000110011001110100001100010000000001110000011000001110110000100111101011111001011011110010111001001000011100011010",
102 => "01001010100001001001001001010101010111101100110100101010100111011000010001110110110111100010010111100101110000001100101001001001101011001001101100010000010010011011110010001100000011101000011010100011010001000000000100111110001000010100110",
103 => "01001110011001110101011101001000011010010011100111100110111110010111001101111000101011000010111111011011111111001111000111000100111100111111000100010101000111010011111010000110000010010000100101111010010111001100100111100100110010010011011",
104 => "11101011010111100100101010000000010001111100010001100100011111011111011010001011110111000010010000010001111101110000000000011101101011111100100100110111111000000000101001111111011001010010010110100010001100011000100001100000010110101010101",
105 => "10100001110001011010100000000111000001011001000001010010001001111001101101101111110011110001100100000111010000110001001000000000001110100011011001010000000001100010011100001100110101100100001011000101110110000001111101111010000010111011110",
106 => "10110100011001101011100101001101111100010011000110010101001000011011100010000110110011000010011100100101001000111000111001001010011111001101000111100011110101111010001100110100100000010001011111100010100100101010110001101000011110110110000",
107 => "01110110111110111100101110110101110001100100100010101010011101010011100000001011010010100011010110000100101010000100100100101111100000101011110100001111110001001001010110011110000110011011010001010110111010101001110001101010010000000000111",
108 => "01011101110100001000010100000100110000101111011111010100111101111111011001011101001001110100110100001100000001010110101000101100010100010001010101100011101110000001000000111111000010011101101110011010011000101110111110100111000100001011000",
109 => "01100110000100010001011100011010011000111111111111111001001010001001111001101001011010100001110111101001000001101110100110111010101110100111001010110111000110000111001000000001100001100000101101110000110110111100110010010011111010100010011",
110 => "01010010100010100111010111111110101000010111111000000110111100111100101001101110111001110001001101001010010110011101111010111011011101010111100101011011000101011001001100111101101110011100011000011000101101011110110010111100011010011010011",
111 => "01001110110001111011110100100111000100100001110100000001110101111111011001010101100001111110111110100011111000001111001000011101001100010110111000011110011001101111101001001100100110111111001110001101001001111101011000000000110000001000100",
112 => "10100101000101111100101111100000010111100111001000110100110100101110000011000100001000011001000000011111110000110101100101110010011100001110110010001010000011110110110110010110010100011100101100000101010000101110100111001011010111001001110",
113 => "00001101010001000011111010011001000110001100001101100000000000011111110000100100111110010011110100011000001100100000100010101010101011010001100010100000111010111011000011101001110001101000110011011110110010101011101101011010101001111000010",
114 => "01101111111100010011110011010011010110110110101000100010000000100000000001110111100110011010011010011001000110001101110111010001000011111001010001011111011011110101000100011110001110111010000101100111101010110110101001110000001010010100011",
115 => "10101111011111111010000000011110101101000000001010001101011110000011111100001100100001000000010101110010111111000100011101001100000011001010100101001000111011101010100101011011010001111111101011001001111111010110001111100011110010000000110",
116 => "00010101010010001001001101000111110111011001010100001101011011111010101100111101100011011100100111100101011011101100000011111100111001001000001110001000101110101011000110100100101001110001110000100110010101101110110001001101100110111000101",
117 => "10000111111001001101111000111010000111100111000100011001000011000110110000100101110010110110111000110110100101111001110110011001010110101110011011010101010000101111011010111001111110100111100111101110110001101001010111100111110110110011101",
118 => "11011001011010100010010110000101001101000101000011010011000001001111101100011100000110101110101100001011110101000110011110110111101111011111100111001101010110001101000011100101101001000010011011101010011111100001001011001000010101011010011",
119 => "10000010110011010001111000000110101100100010011111110110111111111010111010101000101000100101000001110110111000100001100011100111011100111101011000111110101100100011010010000100011011111000000010000100111010001011010001111001011011110010001",
120 => "01100110000011101101100100010101101001000000110001000011001001000100100001001000010101010010110001001010011010100111110001110111000000011100001010011100011001101010010000111110000110011100100011000110001101000010000011100010100100000110111",
121 => "01101000110010101011011010000011101100010111010001111100010000100001001111000101111011100010010100001001010010111011011100101010100101001101001111101111111010100101011000110000010000011011101111010001111111011100001011011110101001111000011",
122 => "11111010111000110101001010000101101110101100000110010010001010111100111010101010101001100000011010100111110001000111100000101100001100111100111011100101000111111110101010010001111111010111011111110010110110010000001111011001001111101100100",
123 => "10110101010101011010101000010001011001001000011010111010010110100101011010110001011111101000100110011100000101110011010001010000001111000110001010100000111100101101000011100011110111000111010110001111110010100001111110100000110000111110110",
124 => "00101101101111110101100010100001010111000000110100010011111011111000110111100100111000110011110111101100101011001001101110011000001111111011010011011100100001000101110010111100110001000110010101011100101000111000000011111011001011110000110",
125 => "10001101011011000001001011111110111110111100001011001000110100001101010111101011011001001110010101110001111011000111101001100111001000011100010010101000101001000110100101101111010001010110101110110001001111000110100100000010001011000011101",
126 => "01011101101100010011011111010100110000000111010000101000111110111010001110000000000100110001001111000001100001011011000011101000010100011001000010001101111101111011100010111110111000111011101000010010001101101101001101110101010010110010111",
127 => "01010000111110000100100101010000010001110001011110101101001100111110011110100111101000001111010111001111111010000001001010000010111110100001111011101111101010001000000111101110101100101111110000011000111111101011001010000110110111001100111",
128 => "00001010110010111010110111000011100110111111101101101100101111101100111000010110001100011110111000001001011101011000110111111110001100010010100011010100010100111111100111010101110011101100110010100110100001010011001100011010100111001001111",
129 => "10001000100011010001000110110111110110101110011100100110101110011110011000010100101010100000101000100000111001100000110110001001101100101101010110000011100010001101110011110000011010110010111000101111001100110010110111001100101111110111111",
130 => "11100111101011010100111100010001000000001001010111011011011110000101101100000011000100100011100111100101100110111001001001101100011001001110011101010111001011111010100110101010111110011000101000110100001100011110111110011101001010001111110",
131 => "00111111011110011110000010100100111010110010010101110000000101001000001110101111001101110100110011110101110010111001000100110011100101101101011010001000100001001010011011100111000110100011010001101001011001110010110011101101000100010011011",
132 => "11111000110010001010100010000101111001001000101010000001011100110011010100010101000100111000111110100010000101110101000010101110100100101111011010110101100011110000111100011101101100111110111111011101111010100011101010110011011010101101111",
133 => "00111110000111101001110110010110100100111111001011000010000101101000001111100001111111111101110110101110000110101111000000101110011111010101000101011001100010111001111110010011001110001110010010111000000000001101111101101111001110000011111",
134 => "00010001010010011101111001110111011110110010011000111100010000000111100100000101100100110010100101010100100101011001111000100101101101111111000010110100010111000111101101010101010111100101111000010110101110000111001101001010101100001001001",
135 => "00011111000101001110001010000101010110111000111010010101101111100110001100011110100010101010011011010001001100000101010010000011010111101001011000101100101010100110011011100100010100011100000000101000100111000110001010001000001101101000010",
136 => "00010110110011101001100001000001101000100001110110011110011111101101100111111111000100111111001110000101000010111010100111001110110011111011011100110100011111001010100110011010011100010110111011011111000111000011001111010011010101101001101",
137 => "00101111000000101100001010000100101110010100101111010101101110100011011110111000010000101000010011111100010111100101101100011010111100111110110111010110110100110111010101010100110111100110000010100110101110101110111110011101011011100010000",
138 => "00111001011111011101100000000111101101001100000101011100011110001010110111000001110000011010011001101010100110111001101111111101001001111111101011001100000010110111100111100010111011000010000010011011001101100010110000110101001010001111101",
139 => "01101011000001001100101001110100001010101101010011001000100101100011011000011011010101011100010000010010011100010011010001111001000010100001100010000110101010111110111110001000000011010110110001111000101001110001111000111101010010010101010",
140 => "00110111010011110010100010101010010011010001001101101000110001010100000110000001110110100100101100000101110111000000000011001101010111010101001100101100110010110100101010111111000110001000110010110111100011010001001000101101110010101100001",
141 => "01011111001111111111001000001100111100111010000011100010111111010101001001110101011111100010010011100101000001000000001010000000101011111101100000001110010111110101100110101110001011110110010000110100111100101001111100111100110101001000110",
142 => "11011101010100011010010010100011001001111111101101010111100010010101101110001001011101110110111000100001101011110010010000001110110001110111111100000011100010010000100100100100101101010000010000011001000110111110101001011010111001111111111",
143 => "01000101101101101111101101001000011110100100001000110010011110110100101000001100101111110111001001000100101001011001001101101111010011000111000010010100111010111101001100110101001010011111111111101111100010110100111101010000001111001100001",
144 => "11111110001110010101011110001110100011110101001001110100000101111110010110100001000111100001000110011101001110000010011010011110001100001101101010110011010001010011101110010000110111010100110000100101000100100001100011000010111100001111100",
145 => "10011011001011010010110011010000101010111001011010011110000011111111000100110101110100101111011001001100100000010100110001010110011011001011011000000001110011010010011101001111011101111111010110101110000011111100101011000011010100110100101",
146 => "10010001001010111010010001101011110010000111100010101010011010010110010011000110011011011100101011010000100011001001010001101100011101101111010011001101100110111110001100100010101011010101011111111010100100000101101010010111000110000110110",
147 => "11010110101011011001001010001101011010101101100000111000110101000111000110111001001010000101100000100010101001111001010111011010000011001101000011001000100111100011011000100101010001001001011110111101101011100101000100000011010111001001101",
148 => "01111001110110111000111001011001000111011101000010110010000011011001010010110000010110101000111011111110101101100101100001100100101100101111001100001011010100000110111011011011011110111111101010010100001010011110001101111100110100110101000",
149 => "00010010001000111001101101010101111000010001100010100100111011111110011000011010011111010001010010000100100000101011000010001011011001110010011010101000001111110001101011010000010110100011111000101111111010100000001110000010000111010010110",
150 => "01100010001001101110111111100000000001000000101001100010110101001001101011000010010111010000100110110111000110001010101100000010011111001011110011111000000110100000101011111100000100010100111111000001101010110010100000110110000000111110000",
151 => "10011000111101010111111101101001001110101111000100111010111100010111111101001101011011110011011001010101001001110001110101110101011010010011011100110010010011000001011011110100110111101100110100010010111110001001011010010000111101110110101",
152 => "10100100110111100011011011001001100011110011100010111100011011011100000101011110100111101110110100001010011010111011111010000101100001110011010110010100111100001101000000001100000111100010110110101001111110011111011110000010110101010100111",
153 => "11010000110010110010011000100110110000100101001101110001000111001100101111000000100100000001111100110001011000110110100100010110001001101101111100101110110001111101001111011101010100110010111101000001111011111010010011000101111011001000001",
154 => "10110101011010000111101011110101111010001101011100010000111111010100000111000001110010010110011101011111000110001110111011101010101111000110011010011000000011010111000101101110111000110011000001100111011100010000010101111001000001010011110",
155 => "00001100100010010110000000101011011011111101010111000100010101110101000010011010010101001011111100100100001111001110110100111011011000001101000100011111000100100111011010111111110110100001000101100111110010000011100001101010000100100000101",
156 => "01111001101010001101000110000011010010001010110001000100011100110000011010111010000100001000010010011101100000010011111111011110110001001111010010110010110010100100011101000001110000001110101101101010000100101101100111101111101000111001111",
157 => "11100101110100000000001101001011011011101010000010001011101001110000111101100010111011100010010110001000111001110010000110100001100100001011010101011110111101001110111010010111101111110010110110010000000111111010101011000001000110011100010",
158 => "10110010001010100001010101011101010100110000000100111010100101101110110100111100000111010111111100001100110111001101111011101001101000111101100011110111000011001110100010011010100001001011000010101101001011001011001000100101000101001011001",
159 => "00000001000000100000101111000011000001110101100011010111111010011111100001110111001111000010110010011100010110001001111111101001000001000010000100111000011111011001100001101101111100011010011100011000000101111001000111001010011010010001010",
160 => "10001111101010001101011111010011010100011100011001110010001100111111011100101000010001011010010010010101010110000011001011001100101110110100110100011010000011111101101010011011101100110001101111110101011100010010111111101011101110100001000",
161 => "00010100011100101101000110111001100010100010010111010100010001001101101110110010011101001110101100101000001101010110111001000101101100100101100000010111010111101001011101001011111100111100110110100111110000101001011010000001110110001001010",
162 => "11000101000110100111000011001111101101111001101001100101011111111010010101010100100001110110111101010010110111001101111100100111011100011010111111110111110100011110100010010010100001101101000100110101000101000101011011011010010100100001011",
163 => "10101010001010000011000001101010011001010010100001100001001101010001110111100010100101010110101011011100010011110110001100100100011010111011001000110100110100111000100101101110100100111100011100110000111110010100001011111001000101111101111",
164 => "01100011101001000110111010000000011010110101101101010001011101110111110011100011001010101110101001000010101001011111111010100001111100011011101100011101000101011100111101000110101000011000011110110101010101101111101101010100101110101000001",
165 => "11000100010011111000001011011101000101010000011101001001011100111000011101011011000011110100100001111010001011001011100001001111110001000011011101001001000101110010010001000001010001111110101100010100010111101100000010110101010100111001001",
166 => "10110000000100101101010011100011100101110100100101001111101010100101011010001111111110111101101011111101111101111001111101110011111111100000000101110100011110001110110100010100010101110111001101111100100010100010011000001101000111110111111",
167 => "11111011010001100111001111101111111001111100010101110011000000011110110010011111100111100011100011100111100010001001001001100000110001001011101000110101010000110011011111110100100010101001001001111111111110010011011101000000110111111000110",
168 => "11111010100110001101110111010100001010110000011000111100001011100010010100101111011111100110111001011010100111100010001001100111111101100110001011011001100010101100110101101001101010100011011110010100010110110000111100110011101110111010001",
169 => "00000001110100101101100110111100010001001001101010010111010111111001110100011001101111001100110000001100010110101011111110011100101000000110111101101010100001110000100010111000101101011101000001010001011011001100101011111001000010100100001",
170 => "00100110110100110010110001100010010110100001001111101010000001001101110110111101010111001010001101011011111011110110001010100001011110100111010110001001001001101011101000000111000000000010111000011110100100111110010101001100110011111101100",
171 => "01001000011001000111010100111110100100111011100100011011011001101010110011000001000010010110100111100010101001000101110111011111101010001000010101011000100110111010111110101110000001010110100100001111010001101100011100010101100010111110011",
172 => "01001001011001100101011010100110100010001111011111010110111111000100010011101111111100001110110100101010100000010010010000000000110000110111000110100000010000010010010010000011000110000001100101111000011101001001101000110010101111011001111",
173 => "10011010101111011001000101000010001001100100110100100011011010010001001110111111101011010111001011011100001001100000001111100001101000011111111111100000011100000001010000101110010101000111100100100010100001111000111101011001010100001001001",
174 => "11011101000011010011111000110010100000010010100100001101011111110011101010001110001000101100110001000110111011111101101111011011000001111111100011101111100001111110010100001111011000110110111111000001000000110110000010011010011001110110111",
175 => "10110111111111110101111111001101111001101001111001101010011010101010011100101100111101010101001010011111011110011001010001100111001110000100001011011001000101110000001010011101111011011100111011101110100111101101010000000010100011100001011",
176 => "00110100010111110010111110101000011100100000100100011111101101111000110111100010100101100001110110101111101100110010101001001100000101101111110001011111001010001111010000011011111101011011111000000110101100000101111101101001001010110000110",
177 => "00111010000011000000110110011011011000110110001101101000110110100010001001001110010001101110111100010000010001010001010000000110111001101011001010001100000011011100010111010100100110000010110011000011111011001100101010110011101111001000010",
178 => "01001100101100111100111100000001011000011101110010100100010011100110101110101001000010101110111011001011001010000110010010001010110001110110110100111100010111010110100011110011111111101000101101111001100011011111101101000100100001001100100",
179 => "10100100000001001000001110011101110111001110100110000100001101110010011110101001010101000000011101011011100100111111101100111010101111111101000100001000000000110100111110001010000010010010011111000001000000101111100101100000101011111101100",
180 => "11001011001100101011001101101111111101011001100110001011000101000000111011111100101110011000001000111010100100101110110100011100001011000000100101111000010001110101101110010101110110100101001000111111101111110010111010011101100100001101111",
181 => "00010110011011101011111001010100011011011010100101110100100111101010100101010110101010010101101110110111010101011001011111011101010010011111101111111011000100011111001100110001111000100011011011000001101101011100100101111001101111010100011",
182 => "00101011100111001110001000001111011111110110000010110001001001100010010000100110010110111101010111001010110010011010000010101100110011000000100101110110101000101111001111101001001100001100111110001100100010001011101111110111111011111111111",
183 => "00101011011000010100000000101000001101101110011100010010110011110100010110000101010011100101001001100100000011011111101101011100001011111000110010001010010011101111011100001000101010110101111010011000001101010111100011101110100100100001111",
184 => "00001000101101001110001010001111101101101101110100000010110011100000011111100011011011110101010101011010000010010010101000011010110001010100110011101000010010011100011000011000000001100010101110110100011010001110001010111110001101000100101",
185 => "00100111001101000001010001001111000110101101100000001100001100001000111111000101110111100011011100001110011011110111111101100111100011011001111010100011001101100101011111000100100101001111001000110101100110000101010010000101000010110011110",
186 => "11100110000111100011001000000001011100001111001000011010111011010010001100110010110101101101111100011010100101110100111011100111100101001011100011010000101111101101101101111001001001000110110011000000001100111110001110010010010011111011001",
187 => "11111110101100101001000010010101100001010001100010001110011000010100011011111000010100001111011001010111110100101101011101110010110000100011111010101111101011011000110101011000001010011101110110110010001100011100010111101101010000001110010",
188 => "11001011111010100000101111011110011011111011100010001101011100001011001110001011100010000000100010011110000010011110110100110101000010101000000111100100000011110110000010100001011000000000111110000101000011010100101001011000111100010110111",
189 => "11001000001111101110100011101000011100100011101101010010001010110110100000101111101011111110110111111001111010101110110101110000101100000100010110000010001100001010000010000001000111101101111100000010000111001000011010001100010101000111010",
190 => "01100100100000000111110000100110001110101101111111110000010000111011001110001011001010111100100000000000110110111000011010010100111001110101100001100010000101000000101011100010001000011100110111000100101101101101111110000111101101001101101",
191 => "00101110111010001100101001100101010000111101101000110011101000010001101110110011000111101011100000001101100100110000110001100110100000011001111011101110100000100010000100001100010011111111101011110101110111000001111100100100010011011000101",
192 => "11111000011001001100100001000110101110001100101110010011000001000110010101001111001000011101100110111100100100110010000001101100110100110000110010110111100100011010010101111101111101010000111100101101000101001111001001110111010100111000110",
193 => "11001101111101011100001000011100101111101111011111111100000000001011011000000010110101101001011011011111101110001011111100000011001110001100001110011110011000101111111101100001010110101110110010101011111011111100111011001100100000100111011",
194 => "01001101011011011000111000111000110011100010000110010111011111110110001001111110101001000011101000010111011111001100101000001100100001111110010010000101100100111111111100001100110010111010100111001010111101011101001010100111011111000101111",
195 => "11111001011110011001011101100001011110110010101111011100011110110011000010110110111101000111100010111101111101010010100101101110001100010010101111001001000100000101100100000011110111011100000010111011110010000101110010000011100011001111110",
196 => "01111110110100001000011011111011010011010111100011000101100101011011111000101000110111000001000000001111000001110010100000110010101001001111001011110111101100011101110101000001010110001000101001100100010001110110100001111011001110111100010",
197 => "01101000011001010110111000011000010110011011110001010111011101101110100110010111111111011010110111101001000000010001000011001000111101110111000000000010101000000101000100010000111010100111111001011100000100100001111111000111001110100001011",
198 => "00111000110101110011000000110100101100111011000111010001011110011011000001010111011100010000010001000101010001010000101000101100110011110110111000111011101111010100010000100001011100010011011100011110101110110011001010111111101001000111000",
199 => "10110001010011110100001011101000101011111011101001110000011010111100010101101101011011011100101110001100101101101110000100111101110100111010011110001010011111100100101010010001110101000011110001111001000010010001011001101110010010010111011",
200 => "01010010111011100110000100001111111011110111001010010100001100101001000011011001000001000000011010010110001001100010101100111000110111110111100110010001101001000000101011011011000111001000000000000100110011101111011001011100010001101100011",
201 => "00101011010000011010001101001110110001101001100001101110000000010100111000001001111010011111010001110011000001000000001001100000100101010010101011000100010100010111100101111100011011001101101101010100001010000111101110010101101000001101011",
202 => "10001110011110101100011110011000001101010001001110011100100101000011101001110011101101010010101001110000010100010111100011100111001110011111001101010001001001111010111110000010101100010100000010111100000111011100101111010000001100011101010",
203 => "01111110111101001001100000100111111010110000011110000000111010000010010110001011001011010101101001110101001011001100110010100111101000110000011100001100011001011111110111011001011101101110001000100111111000111010010110001110101110001000100",
204 => "00111010000110111001000010111011100101111100110001001110110000110010000101101101110111111110100010101010101000111000111010000111010010111000000110110001100110010111001011100010000000110011010011100011001001010111111110110001010110110001011",
205 => "11000010100111110001010011010001011101001010101010100100101010000000101011110101110001001111110111100011001000100101110000010110010101001101010001010100101101011011011111100011100000010101111100001110010010001010011010100001111111110110001",
206 => "00001111111011001101111011010010101110110001110110111000111000011100000001111000110001011111101100110101111101111001101010011111100011111100110100010101111111011110111001111000010000010010110001000100010111110110111101101100001011111100010",
207 => "11011011000011011001110101001011101111110111011110010001001001000100110101000101111101001111011000110011100110100101100000100111100000110000101010000111101000010100110001011101011000100011000001011110001111011111010000000001000111101110101",
208 => "11100001110111100010001111100000101000100011011010101110000000111010101010010010111010010000110000001010011111110000001001010011110100110011111101011100111100011011001100100011000011000000111011110101010001011011001110001001000000110100010",
209 => "00001001100111111010100100011100111001000111100001111001100010111110101101100000001101101111101100110010010011011101010010111100001101011110111110111110010110011100111101010101001001011100001011110011100000011110010010011101110110010110111",
210 => "10110111111101001010100111110010000111011110110010000111111101101001101111000110110001110011000101110010100110010001110000111010110001100011101100000100111101000111001001111100010001001010010101010111000011010110011110100010110100011111110",
211 => "11011000011111000010010001000001010111111101000111010001100111100100011001000010110101001100100000101001000010110101000101100101101111101111100010001010010100111011101010001010101010101010011110110001000000110110111100101011100000011000010",
212 => "10100110100011100111111110101100111101101100011000111111111001000011111000100110111110100100111111000110011011111111011110100000010101111110001110001011001000011000000000010001000111100101011000001001000111010110110101110111001011111001010",
213 => "10100011011000101001011100111000111101011111000100000011100110100010101110101100000011000010001000111111101111101111100011110110100011111110000111101011111101010110110001001111101000000101011100000110110000000001011010001101101011100000011",
214 => "11010101000110010011111010001001101101100111110101011011111111100111010010000101110010100011011101111101111110111010110111000110100000101110101100010110011011101000101101110110011001000000101101001011110100101100110011001001010101010101101",
215 => "00100100001101001001001011000110101011100100110010010111110110110001011011011101101010011010010001010110100000010010011001000101011100010001001011111011101111011111100111000100101011100111111010101110101110010001010110111010010001111001111",
216 => "10110001001010111000011101010100011001100011011100111100011000100100110011001010110110011110110010010110000001010100100001101110011110111010110110100001111000011011111011110001100110101101010101100000001110001011100010010010100111101010001",
217 => "11111110111010001111111101001000000100101001111111111011111110000101000011111010001100110010001001111010000001111000001111011111000110000101000000110101100000010010100000111110111000011110110000011101110011101000100111110011111100110100100",
218 => "00011111000001000100110001010011011110100001001111101110001011010101011110100101001110001010111001001010100111110101100100010000010010011000111100001111110010000001010101111101100110100011010001110000011010011110110001100000000011100011010",
219 => "01101111111001111001000101111100011000010011011000010100001100001110111111111000101011110010110011110101011111110001101101000100100010010111101000010001100001011010000010100010001101011010101110110001101001000100101010110110101011101100100",
220 => "01101111000001101000011100000010111011101010110011000100101011011011010111010010111011000001010100000111110011011101100100110010000111100101111111101011001000001110011010011110101101011101010010101111011100001011011000000101001000000100001",
221 => "11011001010110000001000001001001100110110011110100000101001010111101110110000001010101111100100010100010011110011010001011011001111011011100000001110001101010011000111101100000001000100010111011001010101001100100010100000000011110011010010",
222 => "10110110111101101110111000011111100110000100011011110011000011100000010100011010001011011011001100000010100110111100000100001000001111101011000011001000100010110010101011011010011101010100110000110001010010101110101111101001100000010100011",
223 => "10100110000000011011110000101000010000001100000011101001111001001100101011001100011111111001111101011010001011011011001110001110000011011010001000001011001111100001101001101000011110100011011010001001101010001010101100010101110110110100101",
224 => "00010110001100001110100010001001101001010101111000010100011011010100110000110000101010001100111101100001111011100110101101100001111100001010110011010101100110101100010111100101100111101100000101111101001111000001010001010101000010011010100",
225 => "00010100101111100101111111110111101001000000100101111100001111111001111111010011110001111111010011000110111010110011110110100110001000010010111000101101001011011111000101001100000101001010000000100001100000110111011111110010011000110101000",
226 => "00001101110110100011001011000000100011001001101111100001110010101111010111000010111001101000010100010000100111111100001011101011111011101011000010110010110011000001001010111001000010100111111000001000111011111001100100011001010011111111000",
227 => "00001010000101001110001101110111000000001110010010101001001011000110100110000111001110110010011100101000111001100000100111100010110110110010010001111011101100100100011001000001111001000011100001100001010111110100010100110101111100100011001",
228 => "10101100111001100000011011101010011100111000010001010100101111000111110010110010011111100011000100100000100000110101110001101101000111100011101000110110110101011001000111110011101011000110001011111111110000110110110011111110001100111100001",
229 => "10011000111000111100111001011110100001101110000101110010001110100010111001011101001011000110001000010001101110000110001100111111101010011000011010001001000100010001101010011110101100110110010101101110101000100000000010100011011011111011101",
230 => "11010001001010101111111000101100111000010011110110010010001011001001010101100001000111110000110100111100101001011010111011111110101000111010011100101111111000011000011001010000111001101111111011100010110001010100100110111100011111010010011",
231 => "10110110100011101111110100001010110010110101111111111010110101011101110001101001001100011001011100011110001010101101010010111011010010111101100001001101101100001101010000111111001101011101110011001111011001110110110010101001100111100010011",
232 => "00100010110011101010000001011010010100010111111101100011100000100011110110100101001110010100010110111100010011010010011111100100010101011001011111001111111100010010100101100001010111111110000010011011111001111100110011010010110010010101110",
233 => "00001010010010011110011001000100101001000101101101010101111011100001110111001000010000101110110101000100101000111010100011011101111011010110101111001010111100100000110001100001000010100001101010101101000110000010001110011010111110000000000",
234 => "01001001001101000100101110011100111011010011001011010101010000010110101111100111101100001111011000111000001101011101100011010000100010001000111101001011011010110010111010001110111110001100001010000100000011000110111110100110100111110111001",
235 => "00100110011100010100110101111110011101010000011100111001110110010100111100011110000110010111011010010110000001111001001101011011011011010111110011101001000001100010101100110011111010011100001100100100100010100000010010110000000001000101100",
236 => "11110011010001111000110010001011110010101001110010100111101001011101101000110010101111101101100111111011101001011100011100010100100111100011010000001111011001010001010000110101000011011011001001100101101111010000010001111101001011111010010",
237 => "00000011101000100001011111011001011000010001010100011101110111000100100111000010010000011011000001010010001100001101101001000000110000000111001001001010000011110100011000001000100010010001110100011100011101000101111101000110011100111001101",
238 => "00100011111000111011001110001000001010101011110110100011010110100000111100111100011011111110110111000011001000011000001110010010101110010101100011000101100110100001100110111111110110111001111110001001000000011111100111010111100111110100111"
);

	constant C_data : C_type := (
	000 => "1101110011001001010001101110110111110000101001110110111101010000001100110101101110011110111000110111100011100000100101110011010001101000000000101111000111100110101101111000011100011000001111001101000100100101101111101100011100001111000010000100110111100010",
001 => "1000001000000000110011001100110010111101011101111100100000010000010000010000100011100111100101001011001110011111001000101110001100101000000101111001101001001100001011011001101000101000001111101111110010010101100100100101110000000010001010011001111011011101",
002 => "0100000000101101001000001001011110111001011110000010001110101001110110111000101100111011110011000111100011110100101100001111100000111100011110001000101010101110000110111010000111010011011100111001111101011000101011011101101100001001100110101011010110001111",
003 => "0011111000010101011010001000000100100101001101010011111100110000000101101100110100111110111101100100010000111010000010100011001100011111101011101111110101101010010000111000011111000100000100001001101110011001001100101110011011000111000010001011000101101010",
004 => "0111101011011001010100010111111000001001110011011000101101011100011110011011101010100000111011100010111110001001011100100110111011011101011101101100100100011000100100011001111001101011100111011111111001111011010100000111110000111100011000011010101011000100",
005 => "1011100010101001101100011010111110000110100011100111010101101000001000001111010111111110011101001010110100111101111111001001111000110101110011111001000010110100111001000010001110110100011100110110100000110010001010110111101111101001000100001011000010110011",
006 => "0011111111010000110101010011010101010110101010110101000111101100110101100100001011000111101000011100101110010111001101011010000010110101110111001101011000000010100110011010010101001111011110010000100011111111001011000111101110010001110111110001000101100011",
007 => "0100100110111011001010101011010010010011011110000110101111010011001010111010011101110101111011010100010011001000111111100001111000110011011111110110100000101101101010010100101100001011010010000111000101000011111001101011110000100010001011110000110111111111",
008 => "1010111111100000000010101100011110110110000001010010010011111101101111000001001110111000000110011100111001011011001001010110101111101000100000010001100111011100100010001110010100100010100110110100101010010110111010000101001001101101100001111111110010000111",
009 => "0000010010101111000110000010100111011000001011111111011001101100011101010110100111011101101101000001000111111001011111110111010110011010101010100000100111100100010001010111100110000101000010011111111111110010101101000101011000101100110110110110101101001011",
010 => "1110001101111000000100010111110110111100010111011001111010101011001011001111110111001010101100111100110100110000001101100010111100110000001001011111011100101010110110000001110100101101110111011111010010110010001101011101001011001110001101110101010001010100",
011 => "0111110011111100111011001110001110101001001100000000000110100011101011111111100101110011000111010011000010011100101100000001101100010101001001111000100110000100011000101110010110101010111101000101101000111100111100110000011011110000001100010010010111110010",
012 => "1100011110101010111000111011000100100011111011110010011001110101100110100010010010110001001100010100000010010010000110111100110111111110101011001111100011111010101101001000011111000110001011010011000110101111110110101100010001100011110000010000001001001100",
013 => "0110101101011000111000110000101000110011010011100110001110111000100111001100010100111110100011110011111111100001110101011001110001100101101111010101001110000000000011010001111111010110111001001110011110010111111110010011101001011001101010010011011111010010",
014 => "1011110000010101100111110001110010011100111001110001000010010101001001001101100001001000001101100110000110110011100100101110100010000100110011010010111011000011011001110110100110101100001111000000001110101100110011001001101001101111100011110101110101010111",
015 => "1010001000001111100011101111110000101110110100001011011110010010010001001110001001110111010011101101000101010101101100010011101011110010001011101111110101010000000001000010011110100001000000000111011101001101010000101001000100000100010110101100111001001101",
016 => "1110000001010100100000111001001100111010111000111110100011111110110000010100101111011100010101000000011001111001100111001101000010011111111101110011111000001000110001101100010000111110100101011111100001111011011001011101101110010111110010100111001001111100",
017 => "1101110101010111101001001100100001111010100011001110101000100110100000100110011110001100110001100001010110010010100001001010100100110011011101011000001100111000111010111101100100100011100001111100010110100010000010000110001011010111011100000011011110111010",
018 => "1010110100010110100100111010111011100001110000001101100111011010001010000111110110111110010101001101110001100011011100100101001010011001000011110110001111110000001110010011001010001110101001100000011011000000111110100100001110110011110000111110010011000100",
019 => "1111111001000110111010111100001011111001001000001100011100101011111001100010010000111001001111000110001100100111011011011110111001000110101001011001010110101010111100111101111100001100011100100001001000011111000011110101010101100011000001100001001111001011",
020 => "0001011010111000001100011101001001001111001001100011101111100010101101110011111100100111010101100010010011110001111001011001100110101110101110010100111100100001000010001110001111100100000011111010010000010011011010100110001111000111001110011010010100011001",
021 => "1101010110110111001101101011011010101101010011001111100000010010111011011100000001001100101000000100110100001111011001110100001010100110000000101110101111000010100010101011101111100100010000100011110000100111000111101110101101001111010111011011011100000101",
022 => "0100001010010001101101100100100101011000000010101110111000101100101111100101111110101111001011101011001110010100110011010111011000100011010101011001111111100101100011010000101110111110101010010111110101100010100011111100101001111110011001110000010101110110",
023 => "0100110001100011010000010100000000010001010011001110001111011101000010000111000001011001010000100000100100111111100010101000001111100100000000011000011100001111110000011101010111111000000010000001000011100001111011001101100001010001001101101100100110001101",
024 => "1000011110101101111000001110000101001000010011111110010001011001011011100010111011110000100011000111000010010010111000100110111011011101010010101101001010101001111011111100100111010000100111000000100100101110101010110000000011101000001011100110011101001100",
025 => "1111001111001110011010000101100010110100011000011000111011001100001000111001110101001100000010101001001100100010101010000000011110000010100100010110111110100111101101111010010100001100010011011001100101000111101100011111010001111100110101011100111100011101",
026 => "1101100001010000011001100111100001101111000111101010001101011000011100011000000000001111101110000010010000010011100001000000110001010010000110100010001101110000010100110111101010001001000001110011101100011000101011000001000101011010000100001001110100100101",
027 => "1111101100010011000001001111011000001001111000000100101100011010111001100001111010011111101111101111111000010110011101001001011101100110000100000100110000100010110001001101001001010100000110000110111000101110011001001011001001010100101101010000000000110010",
028 => "1111100100001010101011101011000110110100001111000111000101101100111101100011110110111100010101110011010100100110010101000000010000000000000011011011100110010110011101010101000111011011110011000110110111101001010011100101011110001111101111100000100011010001",
029 => "0101001100100011111001010001111110000011110100101011000110011001111010101001111011101101110111111000101001111011000110111010011001011111011101001001010001100010001001011101100100011110110110111100001011010000010010011001001001010110011100010001111110011011",
030 => "0101111100101101101011000010111101001100001010110101010111001000011010010100100000011000100001101101110001000111001111010100010011000110001010101010000001011101101100110011111001001010110010101000100011011011001000010010101001011101100110011110101101001010",
031 => "1111100001010100111000011101011101111011000010000011011110011111010110001011110010100100011100100001011001110001011010101111100011101011101000100011110110111111111001110000000101111010111100010001100010011101000100100010011011010000000011000000110110000110",
032 => "0101011011000111110110101010110110101011011101111011000001110110010001000000100010101000000110101111000000111010000110011110011011011100111001001110010011100000011000110001101100011000100100001110001111011011110011110000111011100111011010011101001100001001",
033 => "0111000000110110111100111111000000000010001110000101101110110000111101111001000110111101001010000011111110111100101010000001111101011011000011010011010001111110100110010110000111111110001011010011110011010100010111001011100100001011101111011000001000110001",
034 => "1000100100101101110010000010100110101110100111000001001101110110110111000000010000010011100010000010100100100110000100111111010000011010111101110101010100110100001110011000010111101111101011101101001110110111110011111011100011001010011101111000110110001000",
035 => "0001111010000100111010101011111110011010000011100010101011101010011101100100000010101110011000001001001000100001111111110110110011000111011001010000100100000010101001100011000010011011111001101101011000101111001111100110011000001000100100010111111011010010",
036 => "1111100111001011000101000001100011100101011011110100100101010011110111011000011100010010100101011001101100000000111011000010110011010011010110011111100110111100010010001010100000010110010010101111110110010011001100010010111000100001001010110010101011011101",
037 => "1101000110010001011001110011111010101001111011011000100100010100000111101100100101110010100000100001111011010000100111101001100100001000001010101000101010010101001101110100010100011111100110000110100111101101011111111000100011100100011100010011000100011001",
038 => "0000011111011101110010000011101000100011110111101001101111011000101111001001000101101100111100010101001010011101101001010010010111010111100101111101000111010111011010111011010111000011110011110111001111011011100110111110110000001101000010100100010111001010",
039 => "1001000011010010110100110111111001010011101000011110000101000001011000101101111001101010010101110011100111100110001010000100010110010111010011101100110010010011101111111001001001101110000110010001111110111011001101000001010010001011101101010001100011001111",
040 => "0110111011100001101010011010011001110011001100101111010001011100100100101110001101111001111001000101001011001100010010000011010011101101001101100101100100111100101000010101100100111101111010111100011101001100001111000100100100111100000010110011111011111111",
041 => "1001001000010110100010111011110010010010011001000000011010110101101001011100010100101110110001011001101010011110111001100110011011000100011100111011100101110001100010110000110001110011111000111100100010001001011111110000001110010101110000011110110100110100",
042 => "1101000000110000101111100111111011001100110010111000100111101011010010111001001101111110100101111011100100101110101001010100001011010110000001100010000110001100010100000001101001010111001011000111111110000101111001101001110000010110101000111110011110100011",
043 => "1011010111011111010010100010011110100011001011010011011111001101000001001011001100000101011001001010100101101111100011100100001110100100100110101111110111110001001010000111100100101000111111110100111111100011110101101111010010100011111011111010100011001110",
044 => "1011010110001100000101010101000101110010110000100100000111110000111011000010001010010110011110111111101100010111001000001000100010001001110000100011011010001001001110100101011110111100110111111001110101001110011000110100110011100011110010110110011010100110",
045 => "0010000001001000000001100000100011001110001110001010001111111000111110000011111000110111100101000111011010001111000010011101101101110011100100000100000000111000110001011000110100100001100000100100010000011011101010111101111010011011100111111001111100100111",
046 => "1111111101010001110011110010110001111011010011110011011000111011010001011110001001010101010001010101010000001110111100010001010111001111010010111100001001100000101011001110100101000001001001111101000110110101100010001111001010100001111100000111010000000001",
047 => "0101010000101011010101101011101010110110001000001111101110000100111101001110000101110100111010101111011100101101010011010010100111110000111010100000000101110010010011110011111011011101100001101111001000110011000101101110010001100111110101110011101010110101",
048 => "1010111010111110110111101100110101000110111000111110000010000001110000110101101001000111010001111011110100111100000100110011010100101101110101000110110010010101010000000110100000111010000110101111101010110111101100010110101100110011001010100000101100001010",
049 => "1000110010000011001000010110100000001101010110010110110001101101111110011011010001010001010011111011000111001100010000111100010010110100011111101000001001011001111111110010100101000100000001100101111101001000010100100110101101101101111000010110110110001000",
050 => "0001101001110100011110010111000000100100011010101011110101010000000111100111011111011100101101111110001110010100111000010101001111010010000011011011111111000010101100011010010101100110000000110100000101000110110010001110001101110101100110111000001011100111",
051 => "1111101111111111011001101010001111011010111100111011111001101011000101111100011100000001001001100000100001101100100001110111100000110011111000111101100111100011110010011101100010000111001001111111011110100011010110111101001011001111011101000111011011111000",
052 => "0101011000110001110111101000101100010100001011000111001001101001111010110110010000010100011110010110111000010100000111000101011110100010101110000111000110000110000001101011001111001000011110000101000001101010110010101110000101010001000101000100010001010101",
053 => "1101001111010010010100001100111100001111111001001001000001110011110011100111000011101000101000101100010110101010100110010100000111000011111000101100010010011001011000101100101010110100010110000111110011101100101010011011110011001000011011010010100011110111",
054 => "1001100010000110100011000011110010111011111101110000000111100100100100101101110010000110101001011011011101010010001000111011100001100100100001110110101100000111100000110111110110001001101101011010010001001000101011110110001000000111100010100111101111011110",
055 => "1010000000001000111001110110110010000111000000000001111011110011110111101001011001111010011111111100010000100101000111101000100100101001010000100000000001000101001111110101011010001010000010011010111000000001011111110100011100110000111111111011101100010111",
056 => "0111011011101000111000010101011111010001101001000110011111110001000001000110010100111101001111111001001100001011100000010000111011000001010111100001011100100111000000100000100011000101101000010000100000111110011111110100100100101001110111001111011101111010",
057 => "1100000111001100111100001101001011001111001101011101111110011101011000111111110000010111100000000000010110011011100110010101111000101010101011010011011110111001011011000101111101100001101110100011011100011010001010111100000110100001011101100000101000001011",
058 => "0110010101010010100110000111101000101011111100110110111011111011111010000101000010000111000100011111100111111110000110011010101111101001111001010010010110101101101111101001111110010010011111010011011110010111001010101111110111011110010010001011010101000001",
059 => "1110001101001000110101001001111010101001001101110001000010000111101001110000011000101101101110100100001110011011100100010001011111111101111101011001001101111010101111000100101011011100010010000011111010100000001101110101000001001101000101101100010010011001",
060 => "1100001000111010011011111111000100110001111011011000100100111011101101110100101000100100100001000110101110000100000111010011101011100001111001110110110011100001001000101100111101100101101001000011001100010100010101110110111011111110010101110010110010001100",
061 => "1000000110001010110011010010010001100110101110110100101111101111000110100010101110011110001100111111111011011001000011111000100010010101100111001101111011110110011110001111101010111111101000001010110000100001001110100010101111011011010011010100101011111101",
062 => "0100111010010101010101101001011100111101000111011011001001000001101111111010111111010101011000101011010001001011101010010111101110001101110100011100010000011110101011101101001111110111100001100011010110001000111101111000011001100100110000111010000010100010",
063 => "1110011111101011100011100100001100111100000011010100000111111011000000001011101110100101000010101111001111111011010010010010101101001000000011111110110110111101101111010100011010010001001101110011101101001010110000010010110011000001001110001011001010011111",
064 => "1111111001100110001100010010100110110101111111011100010110000111011110111000000110111111101011001100111011101111110010110010111111010100101000001100111011000011111001010111000110000100010010100100111110000010111000000001110101100011000010010101001111100000",
065 => "1010110001000111000110101001000010001110101111011011011011000001011010001111111000100011111101001011100110001011110001101011010111100011100011111111010111110011110010110010100000100001000101001010010101000011010100101111010110111001001111001011100100001100",
066 => "1101100111010101001100110101100011101001111001111101111111110111001100100101000010001101110000001011100110111001110111110000001101001011011100001111010100000011101010011001001101110110001011101111111000111000110011100001100000111100101000010110001110101100",
067 => "1011101001111101111100010101110110000100000101010000010111010111000100100100111010001000011001110010010111111101010100100101010000101010110101100101101100010001110110100110011000000000000010110101101010100000001010110110110001101011110010011000110110011011",
068 => "0100111110000100000100110000011101110101010010110111110000100111001011010111100001100010001011111110010001110110010111111010100010100010101000110000001101000111010110010111001010101100010001010000110001100101111011001001010111011101111111100100010110001011",
069 => "1100010010000111001111000000000110100010111011010000001111110111011011101000110110111100001111011001101010001101010101010011110111001000011100001010110100001110101111111111100110011011110100001100100101010001000110111011111011101111110100101101101010011010",
070 => "0000101101110010010000111110011000011000101011100101001000011011100111111011110001010101111000011000000111001111000110110111001111110101010101110000011101001100110001100000011101111000111110110110100001100100111111010011000101000100001110101110000100000000",
071 => "0100010100100010111010101001100111101011100111001010000010000010010110111101111100100110001010100010000101000000000110100100111100111111111010101101000111100110111101001110010110110101111010111000010100011001011001000011111001110010111101101100000001000001",
072 => "1110010011110101000100101001010101111001000101010011110100111110000100101111010100001010111101000101010010100000100000010111111100010100111010101011101001111000010110110011111010111001110110110001010010010100101001111111110101111000111001011000000110000111",
073 => "1011101011101010001010110110000110010111110001111001000101001000100111111011111111100000000010011100001101001111101000001100110000000100101001000010001111100101001111000001100011001100110100001010001110101111011100011101100101100111011001010011101010111101",
074 => "0000110101000100011100111000010100110001001011100001110110001011101100110010101000101001101110111001011101000110011011010011110100010100110001001101100000001111110110001010110110111010101101010011100100101110010011000111000010001011101010111010001111010100",
075 => "0101001110101011101101111101010110111010001000100111100011010101011110001011011110001110110100100011101100001001001010100001000011001001110101000101110010011011011001010110010000001100001100010011011010100110100000010101101011001100000110100101010100000010",
076 => "1000001111110011000011010110010001001001110001100101001111100111000010111110100010010111000111111110110111011110000110111010010000010001110100110001010110011010100001111110111101111000000111101010100111011010000001011101001100000101010100111010110110010101",
077 => "0101000100101001001011100110010110000110101100001101111100010000000011110001101001111011001010111000101001101011111111100100100111011011100001010110000110000011001000111010111101001111010001001011011100001101001011110010000100010100101100101000100100100101",
078 => "0011000111000000100100111011001000100011100001100111110111010001100110000100001001110100101010101010111011110010001000000010010110110001100100000010011010011101010111111000111011000110101011111111011000110000101110001100101001111000001111000010101110010011",
079 => "0011001100011001100100001001010010001001010001110010011100010000111000100101000110001110001010111000100011011101001011000101010100111110101111101101000100100001000011111111110000110001110011111000011111111101000000110010010001010111101000000010001100100000",
080 => "0111110011001110101101101001010111101001101010010110010100111101010000001110000111011100000000110010111111100011011111010110100101000111001010010100000011100100001100110100110110001100011011000111110001101111101110111001100011100000001010001101111001010111",
081 => "1010110111011011000011010000000010100110001101011101100011110100010001000011111100010111101011100001111011110110010001001101110000000100011111100110111100110100110000101010100101010011111100000101111101001111101110101000110101101000010001111011101111010101",
082 => "1010011101011110010001110100010110100011010000000110001010011110110100101100100111110011101000000010000100001110110000010111110111010100000001110011010100000101010010101100111100001100100001101011011101110001110010010111101110111101101010100010110010001011",
083 => "1001000011000110011101110111100111111100110001110111110100010010100110101100111010000101001110010100101010000000011000101001001010111110100111111100111011011011010100111110100110011010011100010101111000101001010110001110010100011011101110001111011011101110",
084 => "1011000010011101100010101010110111111100110100101000111011111110110000010010010111000101000001101101001111110100011011100101000001000101000011011011111110100111000011111111010000101111110011110000110101011000100011111011101110011110100110101000010110110110",
085 => "1111111110010100111101000010100100011111010100101101111001010110000011101000100001010100010001011010001111101011000110001111010000010100000101111010011110010111111101011110010111010001111001010111110110111111011101000001111101101110000010100000010110001011",
086 => "1000001110111111011100000110010000011111010011100011101000111000110101111001000000100100000111100001101001011111000001110111101001111111110011111100100110000100001011111000001011100011111001110100000000001000011010100101010101111010010010100010010000001001",
087 => "0101000101001101111001000101011110101010101101100101010110110011100010101000100101000100101111010010010001001011111011001000101010011110101100110010011100100010101101100001010100001110100001101000011101111010101000011101011101010011100101101100010010011000",
088 => "0111101110111111101101101011101100101100100000000000111111000100110111001101001000001100001110101011110000000001101010100001010110001101111100000110100010011000110010100110101001101010001101111100010101001111010100011010011111100001011011110111100010100100",
089 => "1001000000101000100000110110101111001111010110000000101001110011001101010111111001001010010001101000010000001001000011110000010110010100100110110111000010100010011111101101111101100111101101101001000101011111010110001000010011000100111110101001001011111011",
090 => "0111001101100010101101100001110000111011110001111111110110100101110100011010101000000000111011011001011110110001011001101100110110100011101001110100000110110111111110011011110001100000010101010011010001101111011001111111001001011100011101110011001011100000",
091 => "0001011010000101101001111001110100100110111010010110100110101000100111111100111101110010000011111011100001010110110000010000101100100100100000011101010101010010000000110000010110000111111100011111100001010111011000100000101101001001001111011111001111110101",
092 => "0010110010100110100000110001010100100001110111111111100000000101100000111110101110010011111101000111010101001101010011101001100011111110000010100011101011010011011111111101101011100100001011111011010100111110110110001011010110000010010010101111010101000111",
093 => "1001101011011100110010001010001101110110010011110011101001111001100100011011001000011101010101011000011110111101011101001110110110011101011101100100110111111111101000001100101011110010111101000100011011000101100010111011100111110011111100100000001101101000",
094 => "1101010011010111100010010111111010011101111111000010000001001100001010011100001011111100100010011100000100100011001001100010001011001001101010110110100101110010011110101010010101111101011100000110000110110011010011100110001110010101001100000110110111110101",
095 => "1111001011110100010101010111010100100011011101111110101010110000001110010011000010101110100110101110011101111111010110100101111100101110100010001000001011110110011000000011100011010110111001001000010100000110011010100000101110111011110010101010110001111011",
096 => "0001011111010011111011011110110100110011101100001001110110011011101010110011101010011001011011011100101100010101001010000011101100111101110001001010111000001101100100110001010110100110000011001101010110001100000010001001010001000000100110100101101100110101",
097 => "0111111000000000010101001011101000100100011110101110111101011001100010110000110010101101000100111100011100000110000110011000111100110011011001010110100100100000001111111011011000110011100101000100011001110100001010110111000111000000010011111010010011110001",
098 => "0111000010101011011001101011100100001101101010000001100011111110101011010001101110001101111111101101101000100101000111010010110001111100011001100001101001010000010001110001100010001101000001001001010001111111011101100101010010011010101010000000010001101111",
099 => "1111000001001000100101110001001000000000100110110110100100001000100001010000001101101100011000011010010110000000111101010001010000010011010100001010101101101001101101101010010101011100101111001111000011110011011001111101000100100111101111010000100000111001",
100 => "0000100000110000011001000111001000001101101101100110100101001110011110011110011101111100110101000000100100001110111000101101100110000100011000001100100010101111010101101110110110111010111011011101110100001000100101100110000100010011101010001001000001100101",
101 => "0100010110110001101100101101110010100001100000100000001100100011010100000100101010101110111110000001101001111000100011010011100100110110110011011100111100111011100100110100011110000101010110011111101110010010000011111001100001000011110100001101011110011111",
102 => "1100101100011010110100101001111101001001111011100100100001110110110001101100110011111001100001100101100101000011100101111010000100001100001100000001101010100000001011011011101110111110111110000110100011001101111011011110111101000001000111111101001010000111",
103 => "0010101100111010011010011001000111111111111110011011100110010111101011100010000100001101111011000110011111100101101010100110011110110001100011101000001101101000100000110010000110110100000101010111111001010111000101100001100010000100000010111100010100111001",
104 => "1010111001100111101001111000101001011000001011000101010111011000101110101101000000110011100111100100111110010001100101110010111101110010001010110111110000001110001010111011101010011010001101111101000100001011001001110010101011111110010010001010001001111100",
105 => "0100000011100101011011101100110100010111000100110001111001101010001111111000100000111000010110100001111111000011100110111110010111010000010110000000000011000111101100100110001101000110010101100011001000100010110010100001110011010000100000010101011011110011",
106 => "0111000001010000111101110100111100101101111000010001011111100011010000000010110000100101000001001001000110110001010110011000110111000001000100111001100111010100010011100011011110100000010001000111000110011110100011100001010111010111011011100001011011100010",
107 => "0001101001101010001110011000111101100010001110011001110100010100110011010101100011101111111100011111000110000010011101100001000010101111011110001000101000110011111000101100000110011100001100111111000100100011101001100011011000100100001001001110000010011001",
108 => "0100000111111001010111111110100101100001001001111111110111011110010101011000100101001010110100100111000100010010001110001100110100110100111010101010001010110011101101011110001100100011110011100110000000010001111111100011111111100101100000000111001100111101",
109 => "1001010001110000100001001000000011011001011011111011111000010100011010001101001101110101010000011001000110001100000111100011111011001010010011110011100100010110011111101011011001000101011000000011101111010010110011001111100110110010101110010010011101110001",
110 => "0011010010100010100011100001100110001111101100100111110110101110111001110011010111111000011001000011000011100100110011011101000001111100111000100001110111000100000100101110011010011000011101111000100110001111100111100111001011111001010100000010001001010110",
111 => "0010000011110000000110001101011101110101100001110111110001011100000011101001100000101111100110101000110011101010100001000101001010111010101100110101000111001100010110100010101111010111111010111001111000101010111110111111111101101010111110111110001101010010",
112 => "0111000000001101010110011000000000110110100110001110100110000001110001101000011100110011101000001111011100100111001011000100101010110110101000010011011010110011001011110100001100011111000111100110000100011010010011100100111100100011011111110100010001010100",
113 => "1100100010111000011101000000110100101101001011010000111111010101011100000111111110000110011001011100101100011111101110101010010000001101010000000100100001110010011110000011001000111001011111000010000100110101010111001010101010101101001011000011000000110101",
114 => "0100110100000101000100001101100110011000000010110110111110000010010110111000100001000101100011010000000100001101000000101111011000000100100100101000011011111100110111001110100010111011110011001101100110100000000011110000010111000110110000000110110010011100",
115 => "0000010001001111111101101001000000010110110110111101110110001011100101011100011001010100101011110101010101000011101001011111111100111111011100010011110110001011101011110101001101010101010100000100010000100111011111000011100101001001001101000101100010010011",
116 => "1010110111010101110101000010111111110100100010110100010010000001011011001111100101101010100111110111011000111110111001011010110011000010111000000100101111111011011011100101001010011001111011010111101010111111001001101011100011011010011001000100101101101011",
117 => "1100010001010110001111000010000010110100010111011010111101000001111011001000001010101011010011001101000000100010001101101101000011000011000100101111000110111011011010100101100101101100011111110100000000011100011010110000000001001011100010000110010010011111",
118 => "1110111101111101011001001101100100001111100010101000011101010101010011001101001001011111111010011111101001101011000100100100110100100010011001011000001010101011111110111110011010010101111100100110001011001010100010010101010110100110100111100001111111011100",
119 => "1000000001111011010001111110010101111100110001011010110001111001011110001000110101101111011011001110100100010100101101100100100011010000111000010001001101011101001100100101011000011101010111000101000110000000000110100111101111010100100110100111000111011010",
120 => "0010001101111010011011000111001111001111111101001010010000111011000111000010000110101010100111100110000100000110011011110000101111001001101011001001010010101111100010000111011000100110001000100000010000111010010011100100010101110011111000111111100110100010",
121 => "1100001000000001000011110101000010000111001101101000101001100100000010001010100111001010100010100011101100100000101110011001011010100000101110010111100100101011110001111001011110000101011101011001010001100000100101111101010010111010111101001010111000011011",
122 => "1111111100111100111010100101010110011110010000001101011010001010011101101100110100100011010110110110110000011110110010111110011010111110001100010010100100110111001110111010010100010010011111011001101111110001011111001000100011111111100000011101100110101011",
123 => "0111000001110110111110001010100101110111101011100101100111000011101101000000111111010001000111110111010010000111101011101001100010010000011100001101000101011000000000100101001000011101100111100000100110000110111001000110110000000111011110110110100101101111",
124 => "0101010110100101001010100111101001000110010111011010110111100111111010101010110000000111001000111001101010111111010111000110101011101100111110111011010000111011100001000101001010111111100000001011011110000010011000001100011100101111010100010011101000010111",
125 => "1010100000011110001101111000110010111010101100010011011000001100111001000011011100010000111101000100000110011001000110111010010010101110101010111110100111001000111101001101000111001111011010111011001100111111010101111101000101001110110010011110111000011011",
126 => "1100110010101101101111001010011000000100100001100001111111010100000101100011100011101000010010010101000000110110110000111100010110011101110000111101011001111000001001101001001101110000111100010101100000111111101001101100100101110111000100100001100000000011",
127 => "1100111111110100101000100110100100000010111110111111110010010110011100101100010000011100001001011110001010010011001001111000010001010011001110010000010110010111011011101011011100000100011010000100000100111011100100010100010010101101010100010100101101110000",
128 => "1101001001100111001011110100101000010001101100101101100011110000100010011010111111100000001000101101011110010100010010100100000101011010110001100000100010101110110011111101110001110010111101111010111111010011101101100001010010110110011011101101110100101001",
129 => "1100111111110111100000110101100010101111001100110010010101111011110110000001001011100111010100011100010100101010100011010000001100100101110010110110011100011000001111111010100001100110100100101000011110001100101010011010010010110001110101000010111101011111",
130 => "1101110110001001100000111001110001100111110101010110111110011110100001000101000101100101001001101100101111100111110010110011110111100110011001001110111101110010111110101111010101011001000001100101110000110000010100011000011011100110010100100110010000010100",
131 => "1101000111011000111110001111000011001110101000101111110010010111000101101011010011110100010001111011100101101111100001110111101111011111010010001010101000100100111010101010000110010000001001001101010111100100110110011100101010011000100010101111110110001111",
132 => "0000101010011011100000000111010111010100000000101100000101101100011101010111111101100000000101001100111011100100011101100001100100000101100111010101001100100000100100100011000100011111010010000100001010101010000101001111111100111101011110110101110000011101",
133 => "1000011110001101001011101100110101101100110010111111010000011100001111100000010001101100111110111000111010100010011110100101100000110111101011110111011011101001000001111000001011111011111000100010111011000110011111000000111100101000110110011100110001000011",
134 => "0100111100001101111010111101110100011100110111111010010100111100111010001001001110100110010110111110100111010100001001010010100101011011111101100010110011000010110100101010101011110001000110101010011110011011101111101000101000111011000010011111101100101000",
135 => "1101101111111011011011001111101101011111011001111001100011110100100100011110101110011010110101000111100110001011011000111010111010000110111011100000010110000010101110000000111000110101110000111011011111111011110011011011010101010111110100111010010100001110",
136 => "0010010101101010010000101001000100101010011101110110011000100110111010011010101111001010101111001001011110110000101111111110111001111011111001001111101001011110001110010001011011010101011010010110100100101110010111101010011110100111101000010111111110001000",
137 => "1111001010100101001001001001111000010001010011101111010100001001001010100101111011110110100100111101010110100111100001111111010001111110011011111011100001111010110000001110111110110100100001100110111010100110010111100101110000000001010101110011100101100110",
138 => "0101011110100011000001110011001100110100001101101010111100100101101001010000001100010111100011001101010101010111100101100001100010101010111000110110111110101101001111011110111011100100001100000011111111100000111111101001001111111010010111001011001100001110",
139 => "1110011010101011101111101101110101010100010101101110111110100100111101011000000011100101100001000011101101111110011000110100101101011111101111111111101111011110010111010010111011010100011100110000110010100100101100010101101000101001100111100110011100000101",
140 => "1100110101110101010111111000001011111010000011101011000010000010110111100001000110101101001101001111011010010011110100100010000110000000011101101000001001000010111010010100011010101111111100111001001011000011111100101011100011001001011100111101010010101000",
141 => "1011001011010100001000011101100010000100101000110110000001101110110100100001100000000111011011101001100001011001101001010010110101111001110000100110011111101100101001000111010010100001110101011010001100010110110000001010100011010110101110011001110111010010",
142 => "0101001001000111010001110101110100111001011010111011010110100101101011101001010011111010100111001001001001000101000011011111000100111001101010101100110101100000001111011100010101000100010100010101101101110001111010110011100101001110111001010011000101111110",
143 => "1111010100100011011100001100101110000111001111101101000101100100100110110100011010011111001001101101001110111010000110100100000001100100110010100000100111010101101011100111110000111110000011000101000110111010111011101010100000000010111000010010001001011000",
144 => "0010000100011010100100010001101110011111111011111000011101110000110000000011111110100101101101011111000000100100110011101111111111011010011100011011011010101010001000001010111101000101111111011111100111001001010111011000101010100100110100100100011111000101",
145 => "0011100000110000111110100010110111011010010011100011000000100100100011100010111111111011111010010011010001101010001101100110100110100100011000000011001000000110001001101101011110001110101010110001100001100100100001010000111010010001111101100110100011100110",
146 => "1010001010100001001101110001011000100100011100000010011110100000010111001110101110111001101010100001110010101100010000010111010100001011100010001000011101001011001100110100111000101110110110111000101000001000010001011100110001111010000100000001001001110100",
147 => "1110101100100010010101110010101110001110100010011100011110000111110101001110011100010111111110011110001111000111001001011000100010101110110000011000001110111111111110111001000110101110001000001100101010101110110000110101010010111000000000000101011111100000",
148 => "1101100001011100011101010011010100001001011111001010001000100110100011101000111100010100110010000101100000010011101110111100111100010101001011000011111001110101100011001111001111111101100100010101001100010000110111010010101101010111111111001001011111111111",
149 => "1111001101010111101111001111010111110001010011111011010000010110010111111100011100001000010110101110000110010101001001111110101110101011111111010010000011010110011110110000001011100010000110011110100001010111111000100110000011001011100010110011110011011111",
150 => "0001011111010100001010100001101001000111001111101111100101000001001010100001111101000101001101010000010010111111101000010100000101100000010101101000100101011110111000000100001010000111010101111100111100000001010111110010100100111010111011011001100000101110",
151 => "0101111010111010001110101100001000010001100101001100110011110000110100100101110000010011110110100110100110111110001001100110001101101100000000101110100000010010011011011010001110000100010100001011101010101011000011011111110111010111101110111000101101100001",
152 => "1100010011011100001001001001011000111101001000110110100011000100111000101111101111000111001001000001100010111000010110010101111101011101010110110111000011001100001100001101001000000010001100011010111010001111101001011111011010111011110000100100001110000011",
153 => "1110011110001001000100100101111010010011010100010111101010011110111000000100011101100010010111101101001010110001011101101101001010000010110011011100100111001101011100110000110000101001100000000100000101010010111101101010000000101010111010001011100010000010",
154 => "0011011100000101010100101111011011001010011010010000011100011010101101101001011001101101111001011100100010001001011110011101011100100001100100010000010010000101000000100010010010000010011101000100111110110111101011111000110101010011111010001101010100100100",
155 => "0000000000000010010100111001000001110101101110010001100100011101011011011001111110010101001000100100100100101110000010110011001010000010110001000011111010010101011111100001010100100100011001101011101101001110111101010000000110011101110000111101110001110001",
156 => "1011110110011110101000010011010011011010110010010110100110000001010001110100111000101110100011000100001100001100111110100110000101101111101111110111011100101011110000101001000011100001101110000000001100001010010000110010011111100000001001100100111010011010",
157 => "0101110110110011100100010111100000001110010011011001110111100001010100111101000000000100011100110010100101110011101100001010111000111010100001001101010101100111110011000110001101101001011110100000001110110110001001110001000101101000000111010011101010100010",
158 => "1000011111011000111110001000100101101010101010100110000010000100100010011110011000000010011110000100000001100001111111011111001010101101011111010011011001011000110101011111001100011011011010010110000100100000000100100000001110010000011101101101001001101110",
159 => "0010011010001000111101010000111001111110111011000101100110010010010110100000010111101010001100000011101100100010111000000010001010101100011111111110010001100001101111010101101101111100100110001010101001111111110111011101011001001110101011001100101110010010",
160 => "1001100001110011100000100011100000111010111100101101011011110111100010111111011011010010101100011010011000110011010111101011001111110100100100010010000011000111111110101011001011000111101101001110100000110110110110111001110011001011000000011111011100111100",
161 => "0100100011111111001001000100110000111110101001100110001101101100001000001001011100101110000100100111110000000101101001100111110011000011011111010010100011111110101010101000001011111111111010000111111101011011011001010000100011010001000001011111001111110101",
162 => "0100001111010010100010100010110111100000000111010101011110101110110111000000011011000101100001101010011101100101110111011010011010110011111100001111100000110110001001110011101010100111000011011110000001111110101101011101101001000000101100000010001110111101",
163 => "1000111001110010100001100101001010011010001011110101111000011001101010111011111111101000010001010000101100011111011011110101101011000110011001011001010111110001110000010010010010001111011000000111110001011100101100011010000101101101000010110010011100011111",
164 => "1000001110000110011000101010110010101110011010001011111000011001011011001000001001011110100010010111001110000001100100000010111011101110101111101000111000000111101110101111000000111000001100100111100111110011010101111100011100000100111100110010111100010001",
165 => "0000000010011000111011001000110001100101000110000000100001101111011101111010001110100110110001111100001101010000100001011100100001011101010100000101100100011100010011111001111011010001110100001110101000110111010001001010110010010011011011010011001100001101",
166 => "1011110100011000000001011110101010100100111000101100111100011010000001011001000100011010001000010000100111100111000001000110000000011111000110011111111101011100110010010011000100011111111000100110000110101110111100101000111100110110001101000010100000111101",
167 => "1110111110010110001001110000100011100101111001110101010010111111111111110110011111010000110111000101100001110010101110000000010110101110111101111110000001101000010110111001001001011111011100011111110001110100110000110010010011001000100100111001110100000111",
168 => "0110110111110100110110100001100101001010010011011111101111010010111001000001010110101011001111100010011100010000110011110011101111110101101111001000111101010110101000010101100101111010010011100000000110111100000100011001101010101100001000100001000011011101",
169 => "1110100000000001001011111101000001100111110010001001010001110111101001011101111001011101011011101100110010000001010100100001010111010011011000000100111101101001010111011000000001100010011100101100100011011111011001111010011111011010110000000100010101100010",
170 => "1010110001000001010010110111101001000101110111011010011111001010110110010011000011011000011000110111100010101010010011101101111101110001001011110011001100110001000100011101010000100110001010101100001001001110101000101111010110101001110110111110001110011001",
171 => "0111010001000000111011111111101100010110001011001100000010101101110101110101110011111111100100011000000010111010101101001110101011001110110010011000111101010110101000110100000111101100101100001000010111010011011010101110101000101111000110111000000100110101",
172 => "1000011110110001111110101101100100011101100110110001100010000010011101101010000001000001010111010110001011011011011101001000111100101000100111000100101011110011110100001101011110010011101100011010000011010011001101000110101101100101001001101101000000000100",
173 => "0010000001101010101010000110110001101011011110101110001111001110000101101001101100010100001110010111001111111011101010111000111110011011010011110101001111110101000110110011011101001000010000011010000001000001011001110110100011000101001010100011011011101011",
174 => "0011111000110000000010100111000101010100000111100111010111100001010100001101010100001010100011100010100110011000101100001001011100110100101011000110100000110110111110000011111010110000000000100001000010101100100101100101101000001101001100100100101010100011",
175 => "1001110110100101010110001111011110100000111100010111000101110010001100111011000010111110101000010011110010001110010101100011010010011110000010010101100001011101110001001010101110101110001011001101101110010101110011001010000010111001110110110110111101111010",
176 => "1010011011101001100100101101010011000010010111111001011101111000000001000111001000000110000100111000110001100111010011100011101110101000011000101010000100111111111110011100000111101101010000001011010100100100000101011110100010011110001101110001011001011000",
177 => "0100110001000100101111110110010101100111011001011101001110000111111011110100101001011111001100011110010011000000110101010111111011100011111000001101110101111001010001100000011110101100000010011111111101010011001000100100001100010010101100101110011111100100",
178 => "1101001101010100011111000100001111111010110111010011110000011101010110101010001010101111000111100111100010000010001011110010001101101100101001110110100000100101110010001100001110100111001110101000011001110001010101110101111100011111001100011100101011001111",
179 => "1100001111101110101011100111100101010101010011011000011011001000010100010110101000110110000001011100110001010011101001001011000100111111110010101100111111010101110100100100110011101010010001001101101110110000000010001011101111000101101000101011010100011100",
180 => "1001001000111100110001101001101101001100000001001110110001101111011101011101101101110001100001001100011100011011001001011011000011110110011111011010110110010100000000011000100101111001000101010111110011000000100110011010000110101000111111111100111001111100",
181 => "0010101011010100111111010111011010111010100110010000111100000011110010111101000000000101110101011001101011000100010110110011110010000010011101101111000110000110001001100101010110100000111001011001000111010000111010110001101011011011100010000001111110010000",
182 => "0100011111010110000111000111000001000011111010100010110010000000111001101100111000101000101000101001001001000101011111010000001111011010010001000100110111110100111101111000001000101101100001010110010000011001000110011010010110100110110000110000111101100111",
183 => "1010011110000011001001101010000110110111000000100100000101111111001000111110101101100010001110010011000110111011101110011110011001101001100101111110101001100101110111100101001110010001000100111011001000101110010000000101101000000101100111111001101000111001",
184 => "1110100010001010111111000111100111110011110100111000110000111001010000101001001011011000000000100001101000011011111100011100001110101101000010010101100100001011011111010100000110100010010101110111100011010000011100001101100011000011101110101000111011111101",
185 => "1000000100001011101110111110111110111100111101010100110110100000010011000010011101101101011100000101010001001011100101001011110110001111110101011110101100001000011101100101011100001011011101110101010001110100010011011100101010101111101100001110101011010000",
186 => "1110000010110110100001111110110110100100111011111110111101110100101011110000100110001000010111010001100010010001001101100111111101011100111101010100110011101111000001101011011011010100111000010110011100011011001100010111010101111110100010001110111010000111",
187 => "0000111110101101001100100111000010010001111000011111000110101101111110001110000000010101111101111101100000111001000111000111001100010010000000010111110000110010101000111100110010001101010101010000011101001101000011011010100100110011010011100001100010101011",
188 => "1110000000000001001010101001100101010100011011011000111000111111000001010001001100111111011001100111110100001100110111001100011111101010100110011000111111001100110001000011111111100011101111111110110101000110100000110101011000110011010001100011101011101011",
189 => "0101010110101111010100101001010000101011111001011001001000111000101110101110010001011010100010100001011010110010010010100011100111011110100111111111011111000101010110001010001111010111001111101100011100001110101111011110111100100111000001110001100101001010",
190 => "0111000111000010010101010101111000101010100110110111101111001100001000000010001000110000101011010101111001101111100100100110011001101010100000010011111001001001100111111010001110111111110011011000111001010100110111110001010100101010011110111110101011111101",
191 => "0000110100011010010011110001001111011010000100000011111010010101011110101111111100100110010101001010110110101101101001000111110000001000000000010111001111011101111111101001111000110010100111101010001001000100001101101001000010000100000101111111110000111100",
192 => "0011100101010000000101111011001111111111100110111111010011111011111000101000100000111001111010010011001011101001010101111111010010001100111010010111101010000110110010001000001101010111101110110111000000101000110100010001110100001011111000100010100010011001",
193 => "1111101111010111010110001100100011100010000000111001110111100100010100000000001100100101101111000101010101110100011101101110100000011000100100010010001001111000100000110100101101110100001000110010110101001011111000101010010010011111000010010100011001111011",
194 => "0001000101010001011101100001101000101001001111010011100000000000111100010010010101111100100000101111101110100100001011100010010011110101010111011111010010111010111110110000110100101000110100011101100100111000110100011011101011011110010110000100101011101111",
195 => "0110100101101101111111011110011110011000111001110011011111100100100000111001101110000011110011110000010100011110010000000110111100101110101111100011100100000101101111111110100000101001110100010001011101100001111100000111001010001000100001001111100100000100",
196 => "1111010110010111010100110111000011111000011101010110010011011101100110000001110110011101110001101000010100001011010101100001100101011101101100110111010010001011000000110011100100101011000000001111011100100101000010110100110110101101110001111010001110011101",
197 => "1011101100110001111100100011010011110000110111110111010010111111010111101100001011001000000101000100010001010001111011011001100011101010110011011101110000110010111011111011000110001010110010111000111011110111101001010100100010001101011111000101001010111101",
198 => "0011101111000001000110001100100110110010010101011100101101000111100110011101001010110011110000010011011110111000011011101011001011000010111010010110010100111000010000010011010111001000000101000111001000011101011001110000110000001111100000010101101111100011",
199 => "0110011110000000101111110110100000110000101110100010110111001110000101001110010100000111001001001101111001000001101100000101010001011000101010111001011011110010111010010101001001111100010010011101000100011000111110100101101111011001110010101111000111010111",
200 => "0111000010110101011010010110101110000110101101111001110101001110010100110101101010011000001000011011000001110110011101010111100110001011010111010011011111010000010100110010010111101110010000110111001010010000010001110101010101101110100110011100001011000001",
201 => "0101110110111000011100000011000110111010010100101001010011011100100111101011001010110010111110101010001101011100110111110111000100011000000001000000010111110000110111011101100001000000100000010111100010010110100001100110101000111011100001011111001111110000",
202 => "1010000100110011000001110011001110010111101110011101110101001000011100110000011010100110100001001000010010011011001100111100111101111010011101000001111111100010100100010100100011001101101100100110001001011001000000011011110110100101100011001011000111100101",
203 => "0011100111101111110111101101110010001000010010101010110000000111111000010011101011111011100110110011100111100110000110101110011101100011111001101010000110101101101111011010100110001101011101111010011000100011000010111000100010010000010011001001101101100111",
204 => "0110100100111101111110101111010101011101111110010011001101001001100010100101010001110100000101110000110101010100011100110111010100001011110010110101111111010110000101111100000101101010110011010101001111100111001010011110001110110000011110000000101000101100",
205 => "1001000111110111010100111011010101000100110010010001010001101000100100111110111111111011111110110011011100000011000111101100011110010001101110000101000001000111001011000101110101101101000011111110100010101011101010000101010010110011101011010100110101011001",
206 => "0110100100110010101100100000110000001111100101100111011100101111101010000101000010100111001011011000100000111101111011100001101101011000011101111101011001001101010011101011011100011000001000100100111010010010000100100100011001111101100100001110101111010101",
207 => "0110000001101000000101100011011001000001011100010101101101111000011011110101011000000110100101000000110010000111001100000110100011110000000110110100101011100101100100011010011000101101001110000110101100111011111110010010000001111011100010110011101101110011",
208 => "1010110010110010011100100110001001100001011010111111100001010010011111000001111111111101110001110001110110111111110011010100101100100100010001100100100111001111010011000111110101110110101101101110000010110101110000101110101100100000100000100111000101011100",
209 => "0010010010011001011000111110100101111100000010100001100011110100011001000000101001111010000001101111010100001111101110000100011000100111010000110111100010001000001111000111001111110101111110101111100011101011011110100011011001011011101001110001000110010011",
210 => "0101110110011100101110010011110001000010101010101000110001110101001000111111111110101010110101111110110000101010111110011000010111111011111000100000101011010110100010110010001000111011101000001000101011011111111110001010101101001001011000100101011100010010",
211 => "0110110001100011100000111011100101100010000110001100000100100011101100101010101100001111111010110100000001010001010001110001001110001110100111001011000110011011011010010000100110110011010000111011011111001001100001011000100011100000000001111110010010100010",
212 => "1010000110000100101111110010100111011010000001100111011111101101101110000001001100000001011111011101000111111110111010000001010001111100011101111110001000011100100010001100110011111111000010110101110001101010000110101111001100101011101001101111000101101010",
213 => "1000111000001111000111110101101101100111000001111000111001110011010001111111100000001011000100001111110001111111000011010001000001110100011101010000000111100000111000111011010110001000010101110101010110011111011111110010110011011001101111001010011111011110",
214 => "1001000110111000000101001011101010110100010110011110100010101010000111110010110110100010100001111111100001001001011100100111001110101111110111110110110110000110111110111101110011101010101011111110011111101110101101000001101101000000011001011011111001111110",
215 => "0001011001001101000101000110111010010101100111000111011110111000100111111111001100000111110100110010111101001000110101000011011011100110110001010001110010101001100010011011010010110110001100110000010001111010101110010100011101110010011001101100000100000111",
216 => "1110001000001101000010100101111101010001100110011101101101101001100001001101010111011010101111011101110100001110100101101111100101111001110000001110010111001101111101000100001001001011111101100111011001111100111001111101001001001111111100111011101110110100",
217 => "1110101001101101001111111010111110011011011110110001010101000100001110001100111110111010011000011011010111110000111111111110101001010110100000111100100001111101101110010110010010110111000110001100110110100010000010100110001011001000100011101101000111101010",
218 => "1111000010110110000111111111101011100100000110000001000000100110000110101010100100000001100100101000001111111010001101011001101000011100001111000000101000111010100101001100100011010111100100011010101100001110001110010111001001011111001110011001111100111100",
219 => "1100101101101110101010111100111110011101011110110001101001101001000101100110111101010111001111000011001001000110011000010110101010101000111101110010101100100000001111001101111001001110101010001000101011101000010010011101000111111010110110101110000100011001",
220 => "0110010011111101111001101101100100100110001100001011010011010110011111101100010011010010001100010011111001110010110010110110100011110111010111100000100000111001101100100110011010001101100111000100101110010010110101110000001000101011010010010011110000100000",
221 => "1101110110111010010001001000011000110001001010101100001010110000001001110111000000001010000100011001101100001010000011000100001101110100011111000010101001001010000011100011000000101011110101111110011111010010010011000001100110011010001011100000110101011111",
222 => "1001111010111111000011011110000011011011011101111000000100011010110100111110110000000001000100110100001001011100110101001100110110001110100000101111011010011001101000001000101101000011101000101011111100010000001110011101000001001100111001111001100100100001",
223 => "0100110010001110101010010101010110111011001100111101011110001111101111101110110101111111110011110110110000001100100111010010101000111100111110000111000001101110110101101101010011001110010100101011111001001101110111100100101110110101000010111000101101001010",
224 => "1011101000110111110000111101100101010100110000011010100001111001101110101011011111011101100101001010100100000101010111001101000111000010000011101000100111001000110010011011100101111111000010100101001001010100011101001101001100010001111000101100000011111010",
225 => "1111100110010001110101111110100011011111110110010110000011111111110010111101010010100111011100111011000110110111100101110001001100001000110111101101100111000001011001010010011000000010001111011010000110001100011000110100010101110110110001001111001001010110",
226 => "0001001010001100101100001010100011100001110111001010011001010101000111001000001101110101101101110011001000100110011000010110110001101111011000111000000101001001100010001000101011010110100010100010111001110110000011000101110001011110010011010110100110010011",
227 => "1110011010111001001110101100000010001110111010001101010010101100110000001001000100101000100000100010100010101000100011101010000111010111100001011111110110010110111111111000110001001101100011101010110000111101011000101100010100011011011001100010111111110100",
228 => "0110111101010010011000001001110101000110001101110011110001110001001111011100000001111110010010101000010111100110101111010010111111101100011110010011010001000101110010111111100111010110011000010011110100011111010011001011010110100111111010100000001001111111",
229 => "1000101000001111101010110010110101110100011100011100001011011111010100001010110111111110111111000100110000000000110000110110110111000001110001110001010111100010000100110010101101110110101001110011001010000111000011111011000000100111001110111110100001100111",
230 => "0000001100101100010101001011101110110100000010100000100101110011000000100001000110001100101101010101110011100100010011010111101001001001110010100100101100011000101111111111001110010011011000001100110010001111100011011111000101111101001011110100011011000001",
231 => "0010100111001110001000000000000000010110011110110111110001010111011101010011000101110110011011001010001101100010011011110101101001010000000100100100111110101101000101111011101010010110011010011000100100101110111110110100011111101110101011100110001110010011",
232 => "1010101100111101100001100001101011100000000001000000100110000010111011100101001001101001011110111111000011001011110010100111000110101011101011111001001001001110010111011011110001111010001100111001100011110011001110011001010010101100000011010000010000001011",
233 => "0110110010011001010001111001111001110011001000000111100001100000101101110111101001100000101110101110001000100000001000001011000101101000001110111110101110000100000100100111001000111110100111100111101111100111111000100101101101101000101100111010001110110001",
234 => "0010000000001111111011100111011100101110101110100011010100101100010001111100011010100011000010010111110111101110000001111001011001110100011000101010011100100010000000101001001000000010011111000101001100000101011000001010010010110111001010001110101001010000",
235 => "1000101010101001100010011100110111111100001010100111101101000101001011000000011100111011010001111110110101001000100001000000010011111110101100101001100000101011111101100010110100011011011001100111011101101000001010110010000001110100101101010111101100010001",
236 => "1111111001110010001100111011111100000011111100001101001011100010110111111100111100110110001101001101101011010001100111001011111111101100101001101111010110111000000100110010101010111011110010111011000000010001011000110101000110000100100101110011100111101100",
237 => "1111110010100110000111011110000110011001101110111111111111010001101110111011100111001101011100101110011101010110111100101101101111111101000101100010010010101101011100110001101111001111010111001111110111101010111111010010011000000011100010100100110001110011",
238 => "1101101000010101110001000001000100110011001100100101001001111000111001001111000111100100111011110001000110010110001011111100011111011110101010110101000111011010001111101101111100001111101010110110010111001101010001111000101100011111001001111000000010100000",
239 => "0001110100110110111010100110000100011111110011010011010100001111001110111101111111111110110010101100010010111110001110010100100111011101001111101011110000100001110111111010000011111111000000001111110101010011000000001000001011011011100001101100101011010010",
240 => "0100011101010111000001011010110101100111100101110001101011001010101001011000100001110101010101011001001001101000010111010010001001100110100110100111011100001011000001001000110100101000101000001011001011111011111100011110010101111000111100110111101001000101",
241 => "1011111100011110111111000101010111111100001111100010111110010101000100101111100100010100010001110110001100101101100111100100000000010011101111101111011111100110001010001011010001100100100111011110011110001010101011001111111000111111000001101101010001100011",
242 => "1010110010010100000100111101100100010001101011010110110011010111111000110110011110001111000010000110000100000100111011111000011011001101000000011111101111000100000000110101110100011101011100101001001010000011010011111001101111100101011111010011110101100100",
243 => "0101100101001010001100111010010010011100100011100000101010001110110110111001101001100101000111001111010100000010100011000110010100110100100110110011001011110100000101101101101110101000100100010001011111001111101110110000110011011001100111000010001000000111",
244 => "1010011101111010110110011100000010010100000011000110011110101010011100111101011011101010111101001101110101010111110111110100110111100101110001000000110100111101001100001011101011110100110111110110110110010001010011110100000100011100101100101101100001100110",
245 => "0100110111100011101100001010100110010011110001111000001110110011111010010110000000010001111010010010101111011010100011011010010011001100000011111011001001101001100011011000010000000011101100101011111011000101101111101110100001011101000011100010000011011011",
246 => "0111010000110111111000110000110101011010001101001101011100010110100111001111010111100001001101110011001010100101000010101110000111101101101010000011101011111100100001011101110100001111100101100110111100101100100111110110111001111001000100101001101100100011",
247 => "1001001100111010000000110110101000011010100000111101011110110101111010101101111101010100000100001000100011001100101101111010111010111101110100100100000110011001010111101000011011000010101001111111001001110010100101101010100011001111010010000101101001100101",
248 => "1111010110010001011011000110000100010111100010010101111111001000111110011110111111000111111111001010100100010011101111010011010100110010101011010011110001101111000000110011100011101000000001001100101001111101001101111110011100010110010010010011100101111101",
249 => "1001111001000101000101011111000010110001110000101010010001011111001001100000010010001111010100001110101001110101000000001101010111100001110110010101011110100101000001011000100111111100101000000111111001000101010011110000000001101000011100000100101101100101",
250 => "1110001011001111010111000100010110101111110111010001101110100011101001000001101000100111011100000000001001011000101000010110000101101101110110101100010100000100000001111010001001001110001001111011000110100010110100100011110001001010100000000111001011111001",
251 => "0100100100000010001110001001011000101001011011000000011010010101101010101111011110011110000101111111001001000011001111000001111100111101110111111100110100000111110001011001001011110100001111110000010001000000010110111011000101101101000011110001110110101101",
252 => "1111010010110001011000011010010010001000010000100111110100100011100101110011111010110011001111010011001101010110110101100000001010011010011111010110011011011100010111000011101001110001101110101010110011100101101010110001100011010100001110111111111111001011",
253 => "0010000010011010111000111011001111110101101110100100000011010101101000111011000110010010010100001100111001001010010001100000000011101000000100010110111001110101101001010100001110010111101100110101101001011100101000100010110001000010100000011010111001101111",
254 => "0011010111111011010100100100110011000011010010000011000010010101101011101000111100010101101010001101100010110100001101100101011100110101110001011011000110110001111101110110011010110100101100101010011100101010111000111000010100111010111010100111010001111101",
255 => "0011110101010000100100001000011111011000000110110011010100010101100110000011101100111110011010000100101100010110000010110101111101111010101111101101101100111101011110101101101111011101110101110000000101110100001000110100001011101001110110101010100010001110"
);
	
	signal X_TB : std_logic_vector(238 downto 0);
	signal C_TB : std_logic_vector(255 downto 0);
	signal ok_cnt : std_logic_vector(7 downto 0);
	signal clk_cnt : integer range 0 to 495;
	signal act : std_logic;
	
begin

	prod_enc : product_encoder port map(ADC_CLK_10, SW(0), X_TB, C_TB);
	
	LEDR <= ok_cnt;
	
	PROC_TOP : process(ADC_CLK_10, SW(0))
	
	begin
		if SW(0) = '1' then
			ok_cnt <= (others => '0');
			clk_cnt <= 0;
		elsif rising_edge(ADC_CLK_10) then
			if KEY(0) = '0' then
				act <= '1';
			end if;
			
			if act = '1' then
				clk_cnt <= clk_cnt + 1;
				if clk_cnt < 239 then
					X_TB <= X_data(clk_cnt);
				end if;
				if clk_cnt > 238 then
					if C_TB = C_data(clk_cnt-239) then
						ok_cnt <= ok_cnt + 1;
					end if;
				end if;
			end if;
		end if;
	end process;

end architecture;