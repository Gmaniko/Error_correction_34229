LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

entity Synch_TB is
end entity;

architecture Synch_TB_arch of Synch_TB is

component Synch is
	port( 
		input  : in std_logic;
		clock  : in std_logic;
		output : out std_logic_vector(254 downto 0)
	);
end component;

signal Clock,bitstream : std_logic;
constant clk_period: time:= 2 ns;
signal test : std_logic_vector(29290 downto 0);
signal indexTest : integer := 0;
signal testhead : integer;
signal result : std_logic_vector(254 downto 0);

--Start Pattern:  0110 0101

begin

-- test <= "0000000000100001000100000000000110010100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101100101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
test <= "00000001100011101011001000001011011110110101000010100001000101010101101011010110111001111110111010110000110001000100100011010100111101011101011111010010110010011010101010000111111101000000101101101000101010110110101100010100011101000001111001100000001101000011010110011011101110000011101101110011101100111110100001000110010101010000010111001011010101011101101000100110000001101010001010000010000100111110000101101000101001001101110101101010111000001101100000111010011110000100011000111101001101111011001110010010110111101100100011101110111010000110101100110111011100000111010111111001001001000110110100001101111000101111011100001110000011100000011010111011011011010110011111100010110000101100011000101010100110000011101000100010010011101100101010000001110110001110111011010110011010000011111111000101001001011011110111101011001100001101011001101110111000001110111110011111110000101100001100001101001111110101110001011011100000001001101111000010111011000000011101011100000000100101010001110110010001011010110000100011010001101100100001101000001010011100111111011111111001101100101110010001011110100111011001101010011000011010110011011101110000011101010001111110101011001110101100111011100011010101001110111010111011100000100111101011101011101100000110111101011001010011110100010111011110101010000010110000110101110001101111101111110111010011100001100111101011010110110101010111111100110110110001001010110000110101100110111011100000111010011010110111001110110110001010100110110000011000101111010101110001010111000100111011100010011111111010001000011011100100010111001011110011010110000011011110111000111101001001100000111001011000010001000000001000011000101110001001100011110110010101010010010001101011001101110111000001110110011111100110000010110000011101001010001000110101010000111011011000000010101101010100111011010001011100001111100110010000011101000000011110110110001110111111111111001111010111001111011011100001011001000101011001101011110111111010100001110011100100000100000011010110011011101110000011101000110000101101101000010011011001101001001000001001011001001010001010011011000111001100101110101100001010000000110001011001110110000001000100111101100101001111000111101000110000010111010100000000101000001100110001000111010000011101000110010111111101110100000110101100110111011100000111011001000111001001010010111100101101011111000000010011001100101110101110011110011110000110010011010100001001100111111001110110001110001110000110000001001110001010011001001101100100100100101110001110010000011101110110101110010011011100111100100110101110110110001101011001101110111000001110100100101000011001110000011001111010011000001100101110010010111100001100011101011110111100000100000011010101100011001111011101111010101001010110110001010110110001001100110101101110101001101101010011010000001110011001000110110010110110111101001110010111110000011010110011011101110000011101100110001011011000011101011110000011000111101000011010101000001010001001010001010011110000010101001011110011111110111110011111010110100010011100011111000011100110011011100000111000110011011011001001011110111111111101100011100100000001110100001101100101110000110101100110111011100000111011110101110101101110000010100000100000100110001010101000111011110001000101101010101010101001001110011001110110101000000111100000111000101110010001100110110100010001001111000110001010100010100111010111010001100010011000010000000110101101110011001101000110110001101011001101110111000001110110011001100010000011011101110100000100111010010011000111000011000001100110010110001101111110000111001101001001110001001000111011111001110101010011101111100000011101101010011010111001111101111111011111000011001110001010101001101111110111011111011111101010100011010110011011101110000011101101100000111101100011110101011100100110111110000000111010000110110000010111000101001011100110110100100101111111000010010011011101001000011011100110000001001011110100010010111011110010010111101000010101101100100000001011010101000100000011111110011101001000000110101100110111011100000111010011111101000110111010010010011010001101010010000001010111001110111000000111011100001000111110101001010111101101111100011101010000010011001101001001001101111010000010010000100000110000000101110101011100010100011110011101001001101101011001010000101011111000001101011001101110111000001110100000100011000101100010000001100010001000001010100001011010110001010101110010100001100110011010000001110000110001100101101000111011011100101101010011100001100001011010111011111000101001110000110001101100101010010001011000110110011010101101000110110000011000011010110011011101110000011101000110101111111100110011110111111100100001101011111011000000010111100000011100101110111011010111110100111011101111111010100010101000110100010100101111001011010110101010101001101100010011000011111110101001001000100010001100100111001110001110000110101001111000110101100110111011100000111010100101001101101000011000111111100011101110001100111110101111001111010101101010101110001010000011110011101111010010010011010001100011100010010101010100110101011101100000001111011111010100011111011111111100110011001001000011101110111010111110001100100011010001101011001101110111000001110111100110111011001100100001101010000110010100100110010111010001111001011100110111000100100110000100001010110001111110101101011011000101000011011101110111101100011010100011100010111101000101001000110110100111000111011011100101001011011101100110100111000001100011010110011011101110000011101010101100100011101011101111111111111010011111010100011111000000010101110100000111001011011111110100001110010110110000010001010010001000110111011111000111110000111111001101011001110010010110010011111011100110101101101100111101110110010100000011101100111101000110101100110111011100000111011111000000110110000010111011001110010011001110110101010101001110111101101011111111000010001001110110110100101011000011100111010010100010010110110110010110001100110011110101111001101001101010100101111010110001000111101101111111100101000001100011001100101010001101011001101110111000001110100000010111101100110111110001001110101011111100010111110111010110011011000011100101100110111100100100101111111111000111010000000100010011010111100111011110111100001111011110011100001010011000010010111010001110000110111010101111001110001010101001101101101100011010110011011101110000011101110010110111100111010001011100010110000110000000101110111101010100011001000000100101010110001010000000100011000110011110100110010110101100111001100001011110111100000110111110011010100111110001001101000000100010010010010010010000010111011011001111101101101000110101100110111011100000111010100001100101000100000010110001101110011010101111101100000010111110110000101011111110001001110010000010101100000011011001000100010000000100001110100011101110000101100001001010001100011011010100011011110100011000001001001100101100110010100100101011001010000001101011001101110111000001110101110100011000001000100110000101001001011001110011001110101011110001110010110111010100111001011111001100011110110010001001110010100110100010010010000101011100100011011010100101111100000010001111101100011011101101100110110100000011010001010011010100110010100011010110011011101110000011101110110010110010010000000001100110000100000011010101011001011001011111010000111001110110111010100010001110001111011000101111111110110011101110101010001001010000111010100000001100000000000000101001100101101001011000101011111001000100111000010010111011111011000110101100110111011100000111011011101001000011100001000110001001011111010101110100010111011010011011111100111111100011100100110010101011101101010000100010111101101001011000001100110110000110010111001110101011000000000001010010011101101110000010010100001000010001111001110010011001000110001101011001101110111000001110110011001000100101000011010100011110001101101100010010001011001010101000001100010000111100111100110110010001101100000110010100100110101100001100000101101001101110010101010010000111000100011010100111000100011111100110111010110010011000001110110000000111110000011010110011011101110000011101110010110001001100110010111101010100100110111111110000010111110110000011001010010111001111000010100100010011110101000110011101001011010011110011111100011100101100000101010111011011100100010010111001111111010100101001101100001110101111011010011110111001111000110101100110111011100000111011110011001110110010100000010110110100111001100111000001010001101111110010110000101101010011000100000100100000011111010011110110101110110001100000100111000000011101101111001010101010000010110011011101010101010011010000011011100111101010111101101110100000010001101011001101110111000001110110101001110101000111001000010110111111101101010001110001100010110010101011101010000000010011101111110110110010011101000000100111001001001100010101100011111000111011010010011101101101111010001100101001000010101010101010100001000001111011001011001011010101100011010110011011101110000011101100111010111110110101010000001011011100101110001000000000001001100111010001000011001100111101101111110000100011000001101000001001000001000010100001010100000000010011010010011100000011111101100000000010110010001000001111010111111001010011011000110011010111000110101100110111011100000111010011101101010001010110001100101110001101111001001100000100101101011001101010011001000101100001101000111000011110111001011010001110001100101110010010001001010111000001101010110110001100011101011110101010000000100101110011101011100100111011101011111010011010001101011001101110111000001110111011110110000101000100110001001100101011110000100000001101111110000000001000111100011010100111110000111111011110110110010110011000111000100111010000000010001100011011011011001010001011111011011010000010101000011101010011010010000001001011101010000111010000011010110011011101110000011101011011110100000110001010001001011100110001111111010010110000000000100000010001000101110010111110011010011111000100110001100011111001001010100010100100111001101001100011101001100111011110101111010011100001000111110000101000011101100101010101010111100100000000110101100110111011100000111010011100000011100110110001111101100100101010111010001111010101111000011110010101000100101000010110110011111000011011000101111111100010011001011111011001010100100010110101011111010101100110000110011100111111110100101100000100101000001100110101101110001010000001101011001101110111000001110100111111100101000011011110010111101111011111010111001000010010000110011000110011011101111010111110110110111111001101110111010100110111100110111011100001110111010101011111000001100010111010101101010010010000100011101111111010001101100110001011010100110001000011010110011011101110000011101011101000100111100110001101111101111110010011110011011010011010110100011110110111110011111000101100000001110110010111100011100111011101010100000100110000011110000001000000011101001101101000111001101101011001011111110100001100111101101010001111101011101111000110101100110111011100000111011110001010010111011100010101011110001110000011000000110110111101011011011011100111000010100110001011001011000101011011101011010001000101000010100000100001000111010110010110111011101010101101010010100111000011100011000100110100001110111000111001011111101010001101011001101110111000001110101010101110011000010100000000000100100111011100111111000101110111101001111000010110111110111101001011000110001101011101100101010001111110101011110010000101001101110000000110110100111011100010011011000001101111000101010010110011100110110110001001111000010000011010110011011101110000011101001000100010010101110101110101100110100010101110110100110000001011111111011000100001111101111111010110010110011111111010100100111110000001101110001110001110011010111000100101011100111100011001001011011111110000000000110011101111101110100011010101010110011000110101100110111011100000111011010100000000010100101010011111101001011011000111100011000101101000000011011010010001001101011100000101001101110000001010001010110101000000110000011100110001000100010111110100000011111000001011010101100111100110101100101010101111100001110110001100011110010001101011001101110111000001110100011101110010000011100101101101110111110011000111000001001010001111111101110100100111011001010111001001100101111011110011010001111101100001111100000001110000010100101001111011000011101011010001001000000000110110110011010000110110100011111111100011110110100011010110011011101110000011101011110110011001111100110111011100010001001100100000111011101100010010011101001101010010011101100001001110101100001010010001110000010010010101001110001011001001001101100101100011001100000101100001111010001100101001101111111111111110011101101100011111110100000110101100110111011100000111011111011100110010110100011101011000010011110000111011010110011100111000101001001011011001111010001110001101011110101110010111110011011110100110110001101011011111110010011111110110000010001010010001001101010010010010010110110110101111010010000101100100011010001101011001101110111000001110111101101101101001100010111000111010001100010111000001111101010101000010001011101001011111101100000111001101100001010001001001100010101101011111010110001101110000101101001010110111000011101010111110011011010100011000010011010011011111111111101111000000101000011010110011011101110000011101010111001001001001110000010000100101101010010001100100101011000100000010001010011011011100110100010001100101111011000110011100101000101101011110001010001010111100101100001100011101001001110101001100001001010110010000000100111101100100100100001011110100100001101011001101110111000001110110000111011110001101100100010011111001000110101000100101111100000001101011111111011010001001100010111100100001001001010001001100000011010111010011110011111101000110100101000001010110100101001010011001110110010000111000010110001100101000111111011100011110100011010110011011101110000011101000111000101111111011100110100000001101111100001100101111110011110110110001111111001001110011111101010110111101001111100110001110001100100011001111000001001111110010111000001110000101101110101011010000000100100110101010110010111111100110000110011110100110000110101100110111011100000111010001011010110011011010001101001101011000111111101111111111100010111011010001111100010100111101010010101011001111110100100110101111100111010000101000010100001111110101100000010001101011100000010010110110010101111010111010010001010101010101100011010111010000001101011001101110111000001110110110101110110010101000110010010101010010010011100001011010111001101101000101000010011010000000010000110100101011010001000101111110001011101111111010010110010101000010110011101101100010100010011100111011011011101110101101110100111100011100101010011001011000011010110011011101110000011101101110001101111101010011100001110010101010101010101001101100010010110110001011010011001110010011010011100000111010100010010010101101110101101110010000100000111111001100001010000011010110000000001011011111010100000011110111101101101101101000100110100111101000110101100110111011100000111011011101101101100011011110110111011010111101111000110011001111011110100011101100010001101010101011000001000100011011111101000001000011101000001010001000110011100111101111111001100100111001011111001110101101100100111000101001010010110110110010111110111011100001101011001101110111000001110110010111110101001001110111010100010001111110000100111011011010011101110010000011000010001110101010011010001010001100001101000001001000111000100011100011101100011001001010000100001101100101001110101110110101111111000000111001010000011000011010100111111000100011010110011011101110000011101100011111101110010100101010110111010100010100001101010101001101000111010101001010100011011010111001111001110011000101011010110111111001111110101010111000001000111011000011001110011011011101110001011100011110110100100100100111001011001101101111010001010011000110101100110111011100000111010110001000011101011010001001111011011101101000111100100010000101011000110111100010010001011100101001110100101010001100001110111011110110101010101110100101101100010011110001111001000100011110100000010101101101001000010000000100100110101000111000010000111100001101011001101110111000001110100010000101000000111011001010001111100001111110001110010100111001001110100000010010100101101001000101110101111011100011010011101111011111000100011110010111010001000110011110111101010101010110010101111000001011101011100100101010101110101111111100001110110000011010110011011101110000011101110111101000011111100011110100000101100110101101000011001111110000011000000111101100001010110000001011111011111111110011110101110110010010000010011101011101011000110000110110111001100011110000001001001101101011011110101100101001000011000110010111011010001000110101100110111011100000111011110100001101010010000111100011011111111000000001001111110111100001011110100000111110111011100010001011110010011101010100011101110100011000100111011001011100010111111111000010011001010001000010111100011010011010011001011001011010010111001100001100000001110001101011001101110111000001110111001110001000011111110101011100100111000000000000101100001001000101011110110101110111101001011011011111111100101101011110011110001101001101000011101100101111101110011110011011111111010001101101110101101011000011000000011000111100000000011011001010011000000011010110011011101110000011101111000011111011101111001001111111100001011011010000111011100111101011110111101001010101101001101001010001001101101011111100101111011111010000101011100011111011011000111011000000111110111111001011001001000001000000000111110111011010001110011010000000011011000110101100110111011100000111010010011001011000110000010000101001111000100010101011011101001010010101001001010100011010000010001111100110011110000101110000110111001000000000101100000000100000111011101101001000011010011010101110111000011000011010011000011101000101001010001100010110101010001101011001101110111000001110111101000100110100100000100111100101010010101000001111010011100000110001010000011011001100101000000100010111011001000101010000010001101011001000001111101111011011000101100011001010100110001100000010011000011101101100100110000011000010111001101011001000010100011010110011011101110000011101110100000001110011101011101101110101110101001110001100000101101010111010010100110010110101111100100111010100000110101101110000100000110001111101110011000011011010110101101111100111000000100011100100110110101101000100101100001001111001001101011110110011101000110101100110111011100000111011010100010011100110110101000000001000111100100110011010001011001101110001100111101011011100010010111111110110000000001011101111111111100111100001111111000001111001101100110101011111101010011011001110001100010110111011111011101000100110010010111100011001110001101011001101110111000001110111011100100100110000110011101110100101101010010110000010010111011011010011101100010000000010110111100101101101111010010001101010101101001111110100110001100110001011111111000100001100101000011110100110001101101001110100010111110010001010000000010100001001100011010110011011101110000011101111001001101001101101100010101000111101110001111010010101001101100010100110011110111101110011000101000001101101101111110111010100111100100011001000111000101000000001100011011110111110010001100110001101000010100001111011110111011010101000001001001000010101000110101100110111011100000111010011001001101101000000000101101110110010011100110011100110000011010011010111101001010001111010100100101010011001010110111011110000010010101100011101011101111000000101111100000101110111011011111011011111110011101110110100111011000001000100001001000100001110001101011001101110111000001110110101011101111110111110000111101100101110101011011110101110000100000000001011101100111100100100110111110001010001110111001000111001110111001101111110001110100001001010011000101101101101111000100110101111010010000000111000011000010110000110010001010111001000011010110011011101110000011101100011110100100000000101010010001000010010100000111010000101101111000100010010000111101111101110010110010011001010110011010111101011011011000101011000111101011010001001001111100101111110100101100011100010101010101001101011111001001111011010100110010001100000110101100110111011100000111010011110110110011110111011010001100100101110100010101110101000011111111011000111100000100011110110100010111000011111011001101000001001001111101000011010000110001011000100001001110001001111110101001101011001110101100111011001100110111111111101111110101011000001101011001101110111000001110100101001000111001110001100001100001100111110011001110101100011100110111000111010100111010100010001011111110011111111010001100001010011001010110101111001101011101110100111101110111100100110000010001100011001011100001011000000011011000110011010000000110111100011010110011011101110000011101011101110111110101101010110010100101101101111111011010110110100101011111001101011100001001010011010110110111111001111000111001101100010101001100101001011110100110101000111010111110101000010110000101010110100010010010100001010011111011101101111011101000101000110101100110111011100000111010111011000010111101001000011111111110000011110100111010111110100111111001010100101011011111110010101011110101011101010000111001010111011110010111010101111010000001100000101100011001000010001001111010111101000111100011110001011001110101111100100101110011100001101011001101110111000001110101001001001010000110100011101011100111000101110000000100011010001111000111100101111001110010100001001100001011011011000110111110001000011111101111001001110010011111011111011110100001000111010000011001010110100101000111110010001110001101111011001000100000100011010110011011101110000011101101001001111100010111011111001100101111001101001100110000000000001100110000111110111110101001001110010110000011010010111010110011111000011110111101010000001010110100000001100000010100110001111100111110001110001001110011011000101000100011011101110101010110000110101100110111011100000111010001000111101010001111000010111111000011010111100010000011100100011010001001010110000001000000010110110011111011111101111100100101011100001011010000111000011001001111100000011011001010000100111000000010011111010000011010011001000011111110111100001010000000001101011001101110111000001110111000100001100000010110011011001011000000010011101010001010010100001101101011110000011101001001000011111011001100101101001100001110111101100101101110101100111011011111001000010001100001111110010011011111001100000110110001011001111000110111000000110101111000011010110011011101110000011101000100110011001001100000100101000011111010111010010111011111111101000110110101101110110110000100001110110000001100110101000010010100000101100011011101111111001000001101111010001111001000110100100100100100000101111010010100100110101010001011010001110011101000110101100110111011100000111010111010001111000000100110010010100001111100010101110001000110100011101100110010110010111101000011100110110110111001001111001011100010100000010110110010110011011000100110001100111111110110111001011011111011100101000011000100101110100011101000111111001101100001101011001101110111000001110100010001101111101111001100110001100110111010111000001001101100001100101110111100111110111011001101000011011000001100000010100111011011111000111000111110001101100100001000001011111011001100101111001000111011101101001111101111111100011101110111101000000001100011010110011011101110000011101101101110100011110111110100000000100101001010100011001100100011011011011010111101111011011010000001000000011000111000010010010100101011011001001111000100000101001100110110001011110011110001111000101110011000101101000111011101111111011100000010110101011010000110101100110111011100000111011110101111101101000100100011110001000101110000001101101101000001001011011011101001000100000110001000011100010010101101010011101010010011000000011110011000001110001100011100010011110110001110100110001011101101011000110101010001101110000011110111011110100110001101011001101110111000001110110100011011100011001100110100100001010010111100110000001110000011110000000011100111100100011011111100110101011100010010001111110100011111101100000100101001011101011100101101100101011001010011011011100111100111000101101110011110111001110010110000111000100100011010110011011101110000011101101111111111100110110100000111110110001101111010111011101110011110110111111000011010111011011000010000111110001011101100010110110100110101011111101001110001000010010101001000111000100010011000110101101101001110000011101000011000110011001111101111011000110000110101100110111011100000111011111111101111110111010100000010100000110010011110010100011011100111000000110000001100100111011000110100010001010000101001010001011010111011110011010000101011100101101000011001010100111000101100010110110010101000110000101111100101000010101100111111000010000001101011001101110111000001110111001000000011100011000000100100011010011000010010100000010110110101100111010001010111100100101101011011101110011110001101111110100010001011100011010100001111111010001001010110110101010111010100000111111001010000111000001101110101010100000011011000001000100011010110011011101110000011101011110001101101000101100011001011010000111000010110100100101101011010101010010011001000111101001100111110101111000010110001010110101000011111101110001010111101001000001110100000101010110100110111101010100101110110000010000101001101001101101001000110010100000110101100110111011100000111011111100110110111000111101001000001001011000011110111100000000110001100110001000101101001011111011100011110101100110010110000101011000111101110101001001100111111001000101011111001010101010111010100001111100001010100101001011011000100000101011100001000010010001101011001101110111000001110100000001000000010011101101001001001010000101111100001111011110001010101001000000011010101110001010100111100010111110000100101001100101010110001011101010101101010001000101101111000101001101101001111101001000001101101001011100000011011011001110101111000111000011010110011011101110000011101001000010001001100001111001010100000110100100000101000000101110110100101011110101011111101111000000100101110100101000100000011101110110111001101011001110010101110110110000111110110011110001010000101001011110100111101111001110011010111111000011000001111101000110101100110111011100000111010101011010111011011011001110100001110000111010101011001011110100101011010011111000101010010111000001011011100111101100101000110011010011111101111010011111010001110100110011000101100010111101010000110000100000010001001110011001011010101111010110001100110100001101011001101110111000001110111101011001001011111000000000111101001000101010101001101001001101000110010111000100100101101010000101010100111000110000010100100001000001101010011001100011100011111000011011001110011111101001111111111110000010100110111000010111001111100001110010000011001000011010110011011101110000011101110101000010110110110101000001011101100100000111101111101111001010111010101010100010001100111001100001001110100110000101101110110101111100101001101111100010101001011000100010110111000100010101111010000010010000100100110011010001101111100001100000110011101000110101100110111011100000111010110000101101010000001011101011101001101001110010011111011100110011101101000101000110100111110000101110000111101100010100101011100110110100110010010111000101011001001111010101100010011101101101001011000100000111110001011110100000011011110101010011011001100001101011001101110111000001110100010011000001111111110000111111101001101011001010001010010111011110111011000101010100111101100000011011100001001011100001111101111001000100100111100011001010101000001101001100001001011111000010011110001000101000100000110011110001101001010000111110100101000011010110011011101110000011101100111010000110101111001000100001011100010110100111000111101100100011110001010101110000110010111011100110101110011010000010100110001001100010100110101000000100010100001110100011011111010010101011101111011001001010010000010111100100000011111001111101010111000110101100110111011100000111011000111101010101100010100110101111100100111101010010011101100100000000110010010100111010100111110000000110001011101110000011001011111100010010001110001010000110010100111101010110110000010111101101001110010111011001111010001101101111110011011110100010001010001101011001101110111000001110101001110110111111010111011000000111001101110000101101010011000111110000110010101100101010100010011110111000100010100010111100111001111000110100000001111011100110000110001100110110111100000011011101000010101100010000110100000110011000000110111111101111000100011010110011011101110000011101000110011010010010000100011101100110100111001001000111100100110101101110100011100001101111100000001000010101010110000101110101000101011000010000001101110101101110010000111000010010100100000011111000111001100000100101011001101010010010011111100011100000000000110101100110111011100000111011000000010101010100110111000100111011011101001000010000101100100111111001001011111001011101010011010110110111001101111000001111001110101011100000011001100101110011000011011011100010100101110011110011111100111101000101100001011111011001010101101100110101111101111110100000101100011110011111111000001011110000101100001001010010011101011001111111011110110010101100111111100001001110011000100101001101111101010000011110101100000001010000101010101011110001111110000100101010100110110101110100101100011110000010101010001010111111100000101111100001000010100110001110011011011001111101101010101001011";
CLOCK_PROGRESS : process
	begin
		Clock<='0';
		wait for clk_period/2;
		Clock<='1';
		wait for clk_period/2;
end process;

inserter : process(Clock)
begin
if (Clock'event and Clock='1') then
	bitstream <= test(indexTest);
	--if indexTest < 29341 then
		indexTest <= indexTest + 1;
	--end if;
end if;
end process;

Synch_instance : Synch
	port map(
		input  => bitstream,
		clock  => Clock,
		output => result
	);


end architecture;


