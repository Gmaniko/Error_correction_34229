LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

entity Decoder is
end entity;

architecture Decoder_arch of Decoder is

signal test : std_logic_vector(254 downto 0);
signal S1result : std_logic_vector(7 downto 0);

component Syndrome1Calc is
	port( 
		R  : in std_logic_vector(254 downto 0); 
		output : out std_logic_vector(7 downto 0)
	);
end component;

begin
	
--test <= "110110011101101001111011111010100001101000110001110110001010101111100010101000100111101101001110100001010101110001011100010111000101000011101101000000001100010010000011100010001110101010011011000011111011011111000010000001001100001011000000101010011000111";
--test <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
--test <= "111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111";
--test <= "110110011101101001111011111010100001101000110001110110001010101111100010101000100111101101001110100001010101110001011100010111000101000011101101000000001100010010000011100010001110101010011011000011111011011111000010000001001100001011000000101010011000111";
test <= "111000110010101000000110100001100100000010000111110110111110000110110010101011100010001110000010010001100000000101101110000101000111010001110100011101010100001011100101101111001000101010001111101010100011011100011000101100001010111110111100101101110011011";

DUT : Syndrome1Calc
	port map(
		R  => test,
		output => S1result
	);

end architecture;
