LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.std_logic_textio.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

LIBRARY STD;
USE STD.textio.all;

entity DecoderBCHE_TB is
end entity;

architecture DecoderBCHE_TB_arch of DecoderBCHE_TB is

component DecoderBCHE is
		port(  
		clock  : in std_logic;
		input  : std_logic_vector(255 downto 0);
		output : out std_logic_vector(255 downto 0)
		);
end component;

--TB clock
signal Clock, ok : std_logic;
constant clk_period: time:=10 ns;
signal result : std_logic_vector(255 downto 0);
signal test, check  : std_logic_vector(255 downto 0);
signal counter, countertest, countercheck  : integer range 1 to 100;

--FOR SINGLE TESTING
type ROM_typeSingle is array (0 to 0) of std_logic_vector(255 downto 0);
constant ROM_SINGLEin : ROM_typeSingle := ( 
0 => "0100000111011100100111100101111110011010110000010111010100010010101011110111000011010110100111110000011001111101000101111110110101000001110111001100101001110000010011000011100010110100111101011101101110101001101110010011110000110101010110101111011100111111"
);
constant ROM_SINGLEout : ROM_typeSingle := ( 
0 => "0100000111011100100111100101111110011010110000010111010100010010101011110111000011010110101111110000011001111101001101111110110101000001110111001100101001110000010011000011100010110100111101011101101110101001101110010011110000110101010110101111011100111111"
);

type ROM_type is array (1 to 100) of std_logic_vector(255 downto 0);
constant ROM_C : ROM_type := ( 1 => "0001010011100001101000100010111010111111110010110001001010110010000011111100111110001000011100011100101010001000110010010001011110100111001101001001001010001011100010110111111001000100011110110101111010011011010010011000100000110010010111110001101111111010",
2 => "0011101000100010010011111101100100001100100111100101001111101011010000101000000111000101111111111111010000111000110000000101000001001100110111110100011101001110101000000111101100001011001110110110000001000000000101110101000111100000101111000110111001100011",
3 => "1000110010110001011110011001111000111111001000000011001001100010011000100110010010000001000001111110111011111000111111011111101101111001001110100011000001110101110101111000110110000110100110101100101101110111001010111110010111010000100111100110001011100100",
4 => "1100001100101000001111111001100000110010000111110100011000111110111101110101000011110001111100100100001111111110111111011111100001100010110101011100110010100100010101011010111000110011110010000100001011111000001010100001100001010000111001110010010011110111",
5 => "0010110000010001101110010010100011111100000010111111111110010001001010111000101111000100000001101010100110110010001111010111010110000110000010011110011110101011011000010100110100110011111110011100110000010011110011101011111000010110010110010110001101110110",
6 => "1011011000000111110101110111010111001010100001010011101010000101110010010101011011100111110001001011111011011100101110000001110100110010010111110111010010111000111001000011101100100100111100101000110001011110100011011011000010100001000110001011011110001110",
7 => "0110001110100110111100111001010001000011010010110101000110111000101011011111001000000010101110000100010111001011110000010001011010101110010111011110110000110000111101011100011010111011001110100101101010001110010101011111111101110111110000101101001111010000",
8 => "0001000000001010000001010110101110000110100010000001111011011011111010101101001001100011011110111101011011110010010100011100110011011011111001100001001111111100101000000110011111001100011011011100000101011011010001111111101110100101000100001100111110000110",
9 => "1100001000110010100100010001110110010110100111000001110011011100111110001011100001101110100111010011011101100011001011010111001001110111010110101110101110010010101110111100110110010111010001000101110111101111000111011011001101000011110000111011110000111011",
10 => "0000110101101110101101111100000000011101101011110001001000101100100111000000110101011010110111000010111101011001101000001010110000010101101101001111110000111110001001110110010010001100001001000111101101010111011001110010001001101101001010101010011110100111",
11 => "0000010101111000110110010000001011010100000110000100000100111001110100011111010011111110000010000010000001000010011101000101010000100110101110100100000010110100011111101110011001001111001010000001110101011100000100111010011111111110110000100011110101101000",
12 => "0001100000011011010101001010110000011111000001111101001010110110010100101101110001001001010110110111100111011010010001110101011111100000000011011101100111010000101110111100100011011110100000000001001000100000111011001001100001100011000100111110100111101110",
13 => "0111110001100001001110110000001010000110000111001111001000011001101010110110010000001100001000010110000011011011100010001000101010011011100111111110011111000001000110100111101011001001110011111111111110010111101111000101010110000110000000001111011000001100",
14 => "0110100000010011100010110111101100011001011000100010001011011000001101001101001100100111111010101111111100000111010110110111111101110100001011011110010010100001101001011111001100010110100111010000001111111001000101100011100110111010110001000111101011110001",
15 => "0000011001110101001010110011000011100011000001011111011010110001011111111110001100100000100011010001001000100011000111110001111111000111111011101111111001101011111110110100111110011101111010111001001010110010100011000011001110000100100011111001111111001011",
16 => "1110000110100101000000000000010001000001110011010101001000100011111111100001011000000000101011001000010010010110010111010110010000000111001110010001011110111100111110100100110101011001101000111100011010011000001000000001110100000011101111111001001011110110",
17 => "1101101100111100111110011010000001011101000011001000110000110101011110101001010100100000011101011010001011110101001110000101101000110001100100000100011100000000001001100100011011010011001111000101011011001101011000100111000111110101010001010011101010001011",
18 => "0010010100011100001000111100010001001100111001101011010000110101010000111101111110011011000000000110010111001000000100101110000000110010100000001000101100001011110010101110001000111011001010010110010000111010101011110010111111011001110111001001110000010111",
19 => "1111110101111101111010001110110001010110110001100000100110010110001010010011110011110011100100110111110110110000001010011111011011110000000111011101100001001110000100011101011111001100110001001111100110110010101010100011010001011110110011110110111110010110",
20 => "1111010101011101101011100001010101111111000110011101101011101011110111010110000110001000000100110100110000001001101000111101111001111000110101100111000000011111001110001001111110100100001001000010100001110111111101100011010001100010000010101010100110100011",
21 => "0000100001010111110000010110001110110100100110101111010001010111010100001011000010111000011101000100001110000101111101101111011011110101111001000010011010001000100111101101011101010001110100000001011100110001001111001100010011011010010000100111110001010110",
22 => "0110101010000100101111100101110011010001000001110001011001111111000101110111001011000110011010111101101001010001101000110111011010111011000100101010011010110001101010111100111100111110001110101010110100110000000111001100101001010001100001001111100011111011",
23 => "1000001110100000110110011111110000111011001111010000100001010000010001110100100100001001110011110110000011111011111001000111001101010011010010100011110111101001110100001100101101110001011110100110110100101101110011111010110001100001010111101100100110111010",
24 => "0000111010111110000010101011111100000100101000001100110001101000111010001111000111001010011010101011001010110110010100011001010001110000101100000000010000011001110011101011010010011111001110000001111001110000100010101010010100011000010010010011100100000100",
25 => "1101101011101101010110111110010110011011001000100010110010100000000000000111110000110001110001011010011001101011100101101100110000011110011010001110111101001010011010011101110110011001111111110011000111010100001001101101110100101000101010001010111110001110",
26 => "0011101000000001100100101100001000001010010101110000000011100010001010111101100110010110110101000000101111001011001010111110000011110110010011101101100000110000111010001100010000000001110110010011010100000110100001010101001010001011100100010100100111000111",
27 => "1000100101100001011110000001101110111000000110101111001111001001011001111010111110011110010111111010000001101111011111100110101101111010000110111110000101111001111001011000110001101100101011011101111010110011001001000101010100011001010011011101111000101111",
28 => "0011101100111111000000011010111110001101000010111000010010010100011110101000000001001011000010101001001001011100101110101011010011111001110011101010011000111111001111111111111100110011111001110011101100001110111001110101001010000001100000111000010001111100",
29 => "0000000010000101001111100000010000101011011001000000100110100010111101011011100010111111000000100000000110001000010011111001111110111011101001111001011100000100010001010110010011110010111010100001100110011100011110001111101010101001000001000001001111000111",
30 => "0110011101111101100010010100001100011010111110010110010000010000010000110011001111101111001110000001000001111100001101011100111011100010101000110101011110001001000000011110010111001011000001000010110000100010010111011000011001100110110001000111101111100100",
31 => "1000111110010011111110000010111110110010010010011011000101100011101001111010001011001010011100001000110011001000110101101100111011111111001110001100101010011001101101001001010101111110110110111100001001111111100011100001110100010101111101001010110010010101",
32 => "0011010111110111010100111111011001010111000001010111011000101000011001101001001100110101101100011110011000100001100101111010010010000110001001001111100000101011100100111011111110100000110110011101010100011101110101011011100100110001110111000101000111011000",
33 => "1101101011111111001000111101110111101010001010101001111111101010111010110101110100111000100111100100010010101000110101100001110011011000000001100110110010111100100010010001100010101100100110010101011110100001101101101110110110011110010001100010100110111111",
34 => "0101101111100111111100111010110111101000011101110100111110110011111110101101111011011011000011111000110111010101111000000011000100101101111111111101111011010010110110011110011111111101111110101110001110111100100011010000011111110111100010100111100110100010",
35 => "1101011111101010001011101001001110000110000111011010000001111010110001010011010111001001001111100011010100011101000000100110001011000100001011001010101011110100101001001111010001111100101100001111101101110100110111110010100000001001110100101110101110110011",
36 => "0100011010110100110000100101010110111110001001100011111011010101010010100101011110110110111111111110001110110110111110001101110100100001101101011010100010000111100011101001100100001001101110000000001000100000111100001101110001110010001110001110010100101110",
37 => "0011110101100001001111110011011111111001001100100010100001001010011100011010000010101110111110000111101100111011001110111110000011101000011100111010111001000001010001011001100101110101100111001001111011001001010111111101010111111100101001101101011101010101",
38 => "1111011001010110001101101011000100000001000101000011001111110100111000110111100011001101010100001000010100100101111010101111011110000010011010011110110111001111110101001110110001010101000101101111111010000011001101100110001101110111011000110000010111111111",
39 => "1111001100111100100001100100111110001011011101111011010010100001111100010011000111101000101001011111101011000001011101111010010110000100110100011000001011111001111100010000111001011010011110000001101011111101100011101011011011100110111010011100010010001110",
40 => "0010010000111001011101110010000011011001110100111100110000010011111111111111101111011011011110010110110001101011100101001001101110110111011010001010001001100110111101010000010011011010100101010011000101101111001100011110100000000011100100101011111111000010",
41 => "0100010000011001100011010101111101010001100100000000101011011000001100011110010110010100110011101110111110000110001110000010001100100011011110110010111001101111000000100111000000101000000100110110110101001100001011110001111110011010010000100001110000101100",
42 => "0001111000100111100110100100000001011011110011111101011100111011001011100000110100100111011111010101101011101101111011010011000101000010000010001110101100100010010010111101100000101010101011001110111001101100110101011111101100111010011101010101010011011001",
43 => "1010000100111110001001001000101111111110000011110110010000011001011000111110000000100101011100000010001010011010101111110001111101111100010110000100111011010000111111010110101110001000010011110110111101110100001011110001001100000111011101110000110010100100",
44 => "1000111111001101001111100001110011101010010000111111010011000100111010111010010011111100100001010000000010011111101011100010000011110101001011001000011001111001010111010101101000101000011000100000110010111101111001001111011100111001000110000000110010111000",
45 => "0101111011111110010000001101101000000101011111010011111000011001110111110111010010111101100010100110110110110001111011010110001000111110011000011100101111111010111110110101111001010010111011110010111011101011010100110101101001000000001001110000010010011011",
46 => "0110010010000000100110011001100010111010100000100101110101011001111000011011000110010101100100101000110100010010001011100111011001110100111111100110010011010111011000100001111101000111100000011100000010000010011010100001000111001011110010110101110001000000",
47 => "1001100110010010111100111100111010000001101011110101000011100000010010000001000101110111111001110010101100001101000010100000110110110100011111101111100100101000111011010111100010110111110010101000001001000111010001101111110101100100111111000110111011110001",
48 => "1111111000100101110100110011011000100010000101100110110101000100011111110010010110000111000110000100001101010010011011000111101011101100101101000111110011001101001011010110001001010010000100000100100000010001001011100000101000111010011011001000110110110001",
49 => "1110011011000010101101000011011011000110001000101110001000011000000000100100100011010101001000011001011001000111001111101000100001100111011001111110011001000001101001000110101111011110010100010011111000100111001101010111011001011110110100100100001011001111",
50 => "0111101100011010001010100110101111110010110000010010110100110111100000011101100000111000001101110110111111111000011000101001101100101100110001010110010010101100010100101100011101010011111000101100110111110100111100001111100110111010001011111101000110111001",
51 => "1001001010110000100000110111110001011001101101001111110100110100101100111101000001111011101001001010001000000011110110000011001001011010111001001001111000010100110001100100100111001011111000100111000110110110011111000110011000101000010001111011111100110111",
52 => "0011111111111100101101010011000000010110010100011101010111101111011001010011111111011011001111010010101001000000100010111000000100111110111001111011010100100000100100000010010010100101111100101100011001101100010011010111001001111100000010011011000001011100",
53 => "0000111000010011000010100101000011100100011011101110001001111111111001011110001010001100010110010010011011000011111001110000100110010110101111010110101111110110110100010011001000010000101010100000111011001001000100101110010001100111000011011101001111101011",
54 => "0100011011101110010010001001101010100001101010001110101001001110100110011011011001000101100011110101000000001011011101111111101011110101010011111111101111101100011110110110011010011110101001010111001001000011011111101111101100010101100111011001001000011100",
55 => "0100100000101010101010000000110010111111001110100010011110110101011011100000001100101100000111011110000100011000011111000000000110100111000100000101001011001100010101110110101110001110111011100100111011101111001010010110110100101000000011111101111000111010",
56 => "1111010100001011011101101010101011100101001010111111011000101110110101010111111010011100011101100111111100000000000110111011111110101011111000011011111001111101100000000000011110011000100111111001011001001101111010001111001001011101101001100110111001010101",
57 => "1001010101000110001001101100100100101010000111110010110110011110001001101000001110110010001010101110000001011000110011011100111010011100011000001011000001110101100010111101000001010010100001110111101011110111110010001110100101011011111000010010100000111000",
58 => "0011000110000001110001000011011111001100110000110100011111100111001000010110010111000110000101011001011001101110000000010100011001011001011111100010101001001100011010111011001110010110001101110001010100001100100111010010000111011100000100101010111000001010",
59 => "1000011101001001100011011000101011110110001011011010001010110111000010101001001001110010110001000001010001010111011001100010010001010001011010111000010000000011011101010111101011101011001010000111101110001101010011000001010110100000000000110011011110011101",
60 => "1111010101101110110110110011011110000110110100011100111111010000111101100101101110111111010001100001101111110111110110000110101100010111111010000110110010010000001011110011111000100111010010100110110010111101011001101011001001111100010000111000001100010011",
61 => "1111110001110001101010001110001000101011111100011111010101110000011000100110000111110100010110100011110100101100001110110011111011001010000100000110000000001010110010100011000011111100001010100111010001100011001010110010000101110011111100001001011101001011",
62 => "1011010100101110000010111110111001010001100000001101010011101000011110110000110100000101101011101000001000101011101111100010101110001000100001000010100110111011011001100111101011110011110010001011010011000010011111110001111010000110010011110101010100111110",
63 => "1100001110000011010101010010010100001110111011110110010001100000101010010111110000110110110111101101001101010000001111110111111010110110001100000011010000000111101110011111000100100110000100001000010010101101010110110101110000111010111001000100100110001111",
64 => "1011110100011000100110110111010110010111011001000000000101010000001100101100001011000110000100111011000000010001110110101010000101001011100101110101101100001001100010010001111111001001011111111001011110010101000100101101101001100000111110110001011001100011",
65 => "1010000111101011110100110010010111101101110100101100000100000001100010110111011111100100000111100111000111101110011010001100011011011010000111110011101110010001011000000110111101111010110001100100000100001110000001000110001000100001110101010001111111110110",
66 => "1100000110110110011111011101110110100011011101000110101010101110011011101110001010111010011100011011100011101011001110101010111010000001011101101111110011000000001001100001111001010101110111001100111101001001101101000011001100110110001110010100000001101101",
67 => "0010000101101000000010110000100011000000101010001000111011110010001001100001111110110011110010010101000000001100000000101000000101001110010001110010111101000000111000011010110110011101000010010101001111100010100110101111000110001010000011101000111001100000",
68 => "0010111111100110111111110101100101010111000001101111000000101110111110111010111001101101110100110110111001100110000101110111011001101111001111101000010011010111111001000101001001010010111100001011000111010010010110000101100111111101111100011111100110100111",
69 => "0100010101110010111100111011011000110101001011010010101001010111100111010001001101110001000000011101011101011110001000011111101111110110100010111100011100101000001000011101011011101110101100110101110001001110010001110011100011110111110111101001111011110111",
70 => "0110100000111011111011000001100111100010010000011101110100100001001010001001101000010100110110011111011110111110110000001000001000011010110010010000100011001011001110100000010000011011111110100011011110110001101000011010011101110101100011010101000110111100",
71 => "0011111111001100110010110010000000011010111011001101110011101111110010001000000101100101101101010111100101110101001111100110101111010110000000011000100100101000111110000001000111111100001000100101110011000111101101100000000101001010111111100110001010010101",
72 => "0111001000101001000001000010111101010000010110000111001111100000011110000011001010011110111000110110001101101100000001010100001001101000001010100010110011000101010101011111101110110011111111111001010010010011101101111110100010101010001101101001100010110010",
73 => "1011110111110001010101110100001000010111110101011001110101011111011000110110001011100101001010010101101011101110111001101001111100000110111001000101100010111100000011001101101001001000011110010100100011000111111000001001101000001000100110011100101011101100",
74 => "1101101011000110001000001010111011010111010001100000111100011110100100100100000100100111011100111111000001010110000110000000101010001100110010100110110001110010001100111110111001101111100111111010111011100001111101110110001111011011110111111100001100110000",
75 => "0000000010010101001100100000001111001100111101011011110000110110101011100111011011100000001010111001011001111011110110101000100001100000111110010011110011100010101101111010111100001110010010111001010111110100111011100101111111100101011111001000001000000000",
76 => "1100101110011101101011001011101111011100101011011101000111100010101110100100011101010110101110110110000100010111000110100010010101010111100001000000100101101111111110110011001011000010010001000010010100001001000010000100010111001011110011010000010000010001",
77 => "1001111110100001101000010010111011001011101000001111111111110000000001110001001000100011000110000100010101001101001110110110000011000011010000111111101001011001110010011100100101110000011100111011001101001101001000011001100010110000100001110000010010011010",
78 => "0110111001001001011011010101110010110001000000010100010100101111110111011000000011001000101011100001100010011000000010011010011101100111010000011100100110101111010110111011010110001011011100001110111110010110010110101110111000110000111011011111111011101111",
79 => "0000000111001110111001100010000001000001010100011100001011111000010001101111100011000010100011101001011000101000110010000110000111000001011100001111110000110010010111101101011101101001010010000101011010011001101111000001001001000110101011010000100101111001",
80 => "0001001100000100110000111101010010010011011110001000100111001111010101010111010011010101111001111100011100100011110011010111010101001010010000010110001110001100101110011110101001000101011001111011101101011111100001110011111000110100000100000001010111011000",
81 => "0001010010001010010110101000011000000010001001101110001101101100101111001011011101111000101011001110100001000100001000101011101011111101011100110110111110011000100010010101010101000000111100100011101011001101000010001101101010111010011001010001100101101010",
82 => "0111110100110001110011001001010110001010000100111100010110010100110101110001110111000010010011011010001000010011010110110111111011110000100010101110110001111100000011101011111010101101110100010011111110101010000101111010100011111010001111000111000001010100",
83 => "1110010111101110100011101100000101001110001111111101001011100111101101101011100001010011010000111101101111110111101001010000111011101111001000111111011000101000001011001010111101111000011111010110010011111110101101000101000100100101111110000010100110100111",
84 => "0011111010100001101001010110110010111011010101100100101001001100111100101101010100111010001110011011011100011000001010000100111010010010100000011101000111000001100011011010111010111000000100100000001101111100010011111000100110100011011101101110010101000111",
85 => "0011100011100010111100100101001101000110001011100000111011000011100111001110010010101110110010001000011101010101111101101000111110110111001100000000100111001000001101110010101110011110011101000101110010001011110011011011101010101001111011101111011001101001",
86 => "0001110011011000011101011001101010010100000011100000011100011010100101001011000011011001110001110011010101010100100110110111011111111011100111010110111111001100001111100110100101011100000010000011000011001010100110111011101111011001000001110111011100101100",
87 => "0101011011100101111010011101001010001000101000101001011101100101001110101001010001100101010100101101000110010011101100100001001100110101010111001001101001011101111100010010001000110011010000000001000010011011000101011000001001110100110000100110010001110101",
88 => "0001010010110101000001011111111000000100000000010101000010111110110000111001000101110011110101000010100111011000010011000011110100110110000100010011000110111101010101100111011100110111111111100101100001100011111000100101101000111100110101111101111110011100",
89 => "1001110011100100010010110110101001110010111001011000010000011100101101110010001011011001100000011111001110001110010100010101000010000100101111100000111100010110111101011001111000011101110000010001001010011100111101011000001001100110110001111110001101110101",
90 => "0010101000010111011001100000000100110010110110010011111001111111110010010101101100000000100111001011111010110101011010010010101011011011010100011011001100100101110010010101110101111011001111010101011010111111001010111001001001100110101011000001100101001001",
91 => "0010111010001010110001000000111001000100011101100010011110000011000010001011111010100000101001111001100001010101111010110001000110010100000010111100111101110010101011011110111001011010011000001010111011000001101111001111101011001111101111100100001000011110",
92 => "1000000110111000110011101010011100001011001100100000001111011010100001001001000110110001000111111011110110100001000100101101110001111010001011100000011110000001110011101011010010101011111101100100010101011100101100011100001011001101101011000011101101011110",
93 => "0011111010000100010010111101111001011111000010111000111111100010000101101100100101101000010110000001001100111011110010100001000101000101000011111100011111111010101000111001110010001100111010001001101001101010101110110000101011010111010101011001010111110100",
94 => "1101011100110100010111101010100101101000000011101000001110000001011000100110010111000001000011100101011110000111100001100000101111000110010100100011100001101001010111001011111100010101001010010100000111101010011111001010111110100111001010000001010110011001",
95 => "1101000011010110110110001101110000000101100110111111001001011101101001100000000010010111101010100010001110100110101000110001101110111111001000011000111100110101111001010010010000100011110101101001001011111001000111100001001101010100010001111100101011101011",
96 => "1100000011110011001111111000001001100111001011111111111101100101010100010111100111100110100110010111101100111100010110111011101110000111001000001110101110010010110001011010110000111011001011000100000000101000000010100100000001101011000101000011011110101100",
97 => "0000111010010000000011110101101011100011111001111010001010110110111101000010100110000101011101101111100111111010000110011000010110101100101111010000011011011011001111010010100000000101110011101101001100111000000101110111000100111000010010010100101100011011",
98 => "0100110111101011110010101101001100001010100101001000101101111001001010010100001101011110000001001101001001111011010111100111010101010010100011110001000000110000101111000011111100001101000101001000100111101111100110000101000101101111110111001110100111000101",
99 => "0011101011010111100110110001100110010101110100110001010110111110110010100010100100101101011110111111011101011000010111111000011111101011001100011101111111000101100100101011011100100001001111000101011011110010110101100010111000101001010100010011001100101011",
100 => "0101000101111111111111111110111100110101010100110111110111001011011111101000010001011001100010010011011010110000011011001010110010011110010001011110001101011110011011101110101110100101000100101010000111111101100101010101110110110110001010000010110110011110"
);


constant ROM_R : ROM_type := ( 1 => "0001010011100001001000100010111010111111110010110001001010110010000011111100111110001000011100011100101010001000110010010001011110100111001101001001001010001011100010110101111001000100011110110101111010011011010010011000100000110010010111110001101111111010",
2 => "0011101000100010010011111101100100001100100111100101001111101011010000101000000111000101111111111011010000111100110000000101000001001100110111110100011101001110101000000111101100001011001110110110000001000000000101110101000111100000101111000110111001100011",
3 => "1000110010110001011110011001111000111111001000000011001001100010011000100110010010000001000001111110111011111000111111011111101101111001001110100011000001110101110101111000110110000110100110101100101101110111011010111110010111010000100111100111001011100100",
4 => "1100001100101000001111111001100000110010000111110100011000111110111101110101000011110001111100100100011111111110111111011111100001100010110101011100110010100100010101011010111000110011110010000100001011111000001010100001100001010000111000110010010011110111",
5 => "0010110000010001101110010010100011111100000010111111111110010001001010111000101111000100000001101010100110110010001111010111010110000110000010011110011110111011011000010100110100110011111110011100110000010011110011101011111000010010010110010110001101110110",
6 => "1011011100000111110101110111010111001010100001010011101010000101110010010101011011100111110001001011111011011100101110001001110100110010010111110111010010111000111001000011101100100100111100101000110001011110100011011011000010100001000110001011011110001110",
7 => "0110001110100110111100111001010001000011010010110101000110111000101011011111001000000010101110000100011111001011110000010001011010101010010111011110110000110000111101011100011010111011001110100101101010001110010101011111111101110111110000101101001111010000",
8 => "0001000000001010000001010110101110000110100010100001111011011011111010101101001001100011011110111101011011110010010100011100110011011011111001100001001111111100101000000110011111001100011011011110000101011011010001111111101110100101000100001100111110000110",
9 => "1100001000110010100100010001010110010110100111000001110011011100111110001011100001101110100111010011011101100011001011010111001001110111010110101110101110010110101110111100110110010111010001000101110111101111000111011011001101000011110000111011110000111011",
10 => "0000110101101110101101111100000000011101101011110001001000101100100111000000110101011010110111000010111101011001101000001010110000010101100101001111110000111110001001110110010010001100001001000111101101010111011001110010001001101101001010101010011110100110",
11 => "0000010101111000110110010000001011010100000110000110000100111001110100011111010011111110000010000010000001000010011101000101010000100110101110100100000010110100011111101110011001001111001010000001110101011100000100111010011111111110110000100011110001101000",
12 => "0001100000011011011101001010110000011111000001111101001010110110010100101101110001001001010110110111100111011010010001110101011111100000000011011101100111010000101110111100100011011110100000000001001000100000111011001001100001100011000100111110100011101110",
13 => "0111110001100001001110110000001010000110000111001111001000011001101010110110010000001100101000010110000011011011100010001000101010011011100111111110011111000001000110100111101011001001110111111111111110010111101111000101010110000110000000001111011000001100",
14 => "0110100000010011100010110111101100011001011000100010001011011000001101001101001100100111111010101111111100000111010110010111111101110100001011011110010010100001101001011111001100010110100111010000001111111001000101100011000110111010110001000111101011110001",
15 => "0010011001110101001010110011000011100011000001011111011010110001011111111110001100100000100011010001001000100011000111110001011111000111111011101111111001101011111110110100111110011101111010111001001010110010100011000011001110000100100011111001111111001011",
16 => "1110000110100101000000000000010001000001110011010101001000100011111111100001011000000000101011001000010010010110010111010110010000000111001110010001010110111100111110100100110101011001101000111000011010011000001000000001110100000011101111111001001011110110",
17 => "1101101100111100111110011010000001011101000011001010110000110101011110101001010100100000011101011010001011110101001110000101101000110001100100000100011100000000001000100100011011010011001111000101011011001101011000100111000111110101010001010011101010001011",
18 => "0010010100011100001000111100010001001100111001101011010000100101010000111101111110011111000000000110010111001000000100101110000000110010100000001000101100001011110010101110001000111011001010010110010000111010101011110010111111011001110111001001110000010111",
19 => "1111110101111101111010001110110001010110110001100000100110010110001010010011110011110011100100110111110110110000001010011111011011110000000111011101100001001110000100011101011111001100110000001111100110110010101010100011010001011110110011110010111110010110",
20 => "1111010101011101101011100001010101111111000110011101101011101011110111010110000110001000000100110100110000001001101000111101101001111000110101100111000000011111001110001001111110100100001001000010100001110111111101100011000001100010000010101010100110100011",
21 => "0000100001010111110000010110001110110100100111101111010001010111010100001011000010111000011101000100001110000101111101101111011011110101111001000010011010001000100111101101011101010001110100000001011100110001001111001100011011011010010000100111110001010110",
22 => "0110101010000100101111100101110011010001000001110001011001111111000101110111001011000110011010111101101001010001101000110111011010111011000100101010011010110001101011111100111101111110001110101010110100110000000111001100101001010001100001001111100011111011",
23 => "1000001110110000110110011111110000111011001111010010100001010000010001110100100100001001110011110110000011111011111001000111001101010011010010100011110111101001110100001100101101110001011110100110110100101101110011111010110001100001010111101100100110111010",
24 => "0001110010111110000010101011111100000100101000001100110001101000111010001111000111001010011010101011001010110110010100011001010001110000101100000000010000011001110011101011010010011111001110000001111001110000100010101010010100011000010010010011100100000100",
25 => "1101101011101101010110111110010110011011001001100010110010100000000000000111110000110001110001001010011001101011100101101100110000011110011010001110111101001010011010011101110110011001111111110011000111010100001001101101110100101000101010001010111110001110",
26 => "0011101000000001100100101100001000001010010101110000000011100010001010110101100110010110110101000000101111001011001010111110000111110110010011101101100000110000111010001100010000000001110110010011010100000110100001010101001010001011100100010100100111000111",
27 => "1000100101100001011110000001101110111000000110101111001111001001011000111010111110011110010111111010000001101111011111100110101101111010000110110110000101111001111001011000110001101100101011011101111010110011001001000101010100011001010011011101111000101111",
28 => "0011101100111111000000011010111110001101000010111000010010010100011110101000000101001011000010101001001001011100101110101011010011111001110011101010011100111111001111111111111100110011111001110011101100001110111001110101001010000001100000111000010001111100",
29 => "0000000010000101001111100000010000101011011001000000100110100010111101011011100010111111000000100000000110001000010011111001111110111011101001111001011100000100010001010110010011110010111010100001100110011100011010001111101010101001000001000001001110000111",
30 => "0110011101111101100010010100001100011010111110010110010000010000010000110011001111101111001110000001000001111100001101011100111011100010101000110101011110001001001000011010010111001011000001000010110000100010010111011000011001100110110001000111101111100100",
31 => "1000111110010011111110000010111110110010010010011011000101100011101001111010001011001010011100001000110011001000110101101100111011011111001110001100101010011011101101001001010101111110110110111100001001111111100011100001110100010101111101001010110010010101",
32 => "0011010111110111010100111111011001010111000001010111011000101000011001101001001100110101001100011110011000000001100101111010010010000110001001001111100000101011100100111011111110100000110110011101010100011101110101011011100100110001110111000101000111011000",
33 => "1101101011111111001000111101110111101010001010101001111111101010111010110101110100111000100111100100010010101000110101100001110011011000000001100110110010111000100010010001100000101100100110010101011110100001101101101110110110011110010001100010100110111111",
34 => "0101101111100111111100111010110111101000011101110100111110110011111110101101111011011011000011111000110111010101111000000011000100101101011111111101111011010010110110011111011111111101111110101110001110111100100011010000011111110111100010100111100110100010",
35 => "1101011111101011001011101001001110000110000111011010000001111010110001010011010111001001001111100011010100011101000000100110001011000100001011001010101011110101101001001111010001111100101100001111101101110100110111110010100000001001110100101110101110110011",
36 => "0100011010110100110000100101010110111110000001100011111011010101010010100101011110110110111111111110001110110110111110001101110100100000101101011010100010000111100011101001100100001001101110000000001000100000111100001101110001110010001110001110010100101110",
37 => "0011110101100001001111110011011111111001001100101010100001001010011100011010000010101110111110000111101100111011001110111110000011101000011100111010111001000001010001111001100101110101100111001001111011001001010111111101010111111100101001101101011101010101",
38 => "1111011001010110000101101011000100000001000101000011001111110100111000110111100011001101010100001000010100100101111010101111011110000010011110011110110111001111110101001110110001010101000101101111111010000011001101100110001101110111011000110000010111111111",
39 => "1111001100111100100001100100111110001011011101111011010010100001111100010011000111101000101001011111101011000001011101111010010110000100110100011000001011111001101100010000111001011010011110000001101011111101100011101011011011100111111010011100010010001110",
40 => "0010010000111001011101110010000011011001110100111100110000010011111111111111101111011011011110010110110001101011100101001001001110110111011010001010001001100110111101010000010011011010100101010011000101101111001100011110100000000011100100101011111101000010",
41 => "0100010000011001100011010101111101010001100100000000101011011000001100011110010110010100110011101110111110000110001110000010001100100011011110110010101001101111000000100111000000101000000100100110110101001100001011110001111110011010010000100001110000101100",
42 => "0001111000100111100110100100000001011011110011111101011100111011001011100000110100100111011111010101101011101101111011010011000101000010000010001111101100100110010010111101100000101010101011001110111001101100110101011111101100111010011101010101010011011001",
43 => "1010000100111110001001101000101111111110000011110110010000011001011000111110000000100101011100000010001010011010101111110001111101111100010110000100111011010000111111010010101110001000010011110110111101110100001011110001001100000111011101110000110010100100",
44 => "1000111111001101001111100101110011101010010000111111010011000100111010111010010011111100100001010000000010011111101011100010100011110101001011001000011001111001010111010101101000101000011000100000110010111101111001001111011100111001000110000000110010111000",
45 => "0101111011111010010000001101101000000101011111010011111000011001110111110111010010111101100010100110110110110001111011010110001000111110011000011100101111111010111110110101111001010010111011010010111011101011010100110101101001000000001001110000010010011011",
46 => "0110110011000000100110011001100010111010100000100101110101011001111000011011000110010101100100101000110100010010001011100111011001110100111111100110010011010111011000100001111101000111100000011100000010000010011010100001000111001011110010110101110001000000",
47 => "1001100110010010111100111100111010000001101011110101000011100000010010000001000101110111111001110010101100001101000010100000110110100100011111101111100100101000111011010111100010110111110010101000001001000111010001101101110101100100111111000110111011110001",
48 => "1111111000101101110100110011011000100010000101100110110101000100011111110010010110000111000110000100001101010010011011000111101011101100101101000111110011001101001011010110001001010000000100000100100000010001001011100000101000111010011011001000110110110001",
49 => "1110011011000010101101000011011011001110001000101110001000011000000000100100100011010101001000011001011001000111001111101000100001100111011001111110011001000001101001000110100111011110010100010011111000100111001101010111011001011110110100100100001011001111",
50 => "0111101100011010001010100110101111110010110000010010110100110111100100011101100000111000001101110110111111111000011000101001101100101100110001010110010010101100010100101100011101010011101000101100110111110100111100001111100110111010001011111101000110111001",
51 => "1001001010110000100000110111110001111001101101001111110100110100101100111101000001111011101001001010001000000011110110000011001001011010111001001001111000010100110001100100100111001011111000100111000110110110011111000110011000101000010001111011111100110101",
52 => "0011111111111100100101010011000000010110010100011101010111101111011001010011111111011011001111010010101001000000101010111000000100111110111001111011010100100000100100000010010010100101111100101100011001101100010011010111001001111100000010011011000001011100",
53 => "0000111000010011000010100101000011100100011011101110001001111111111001011110001010101100010110010010011011000011111001110000100110010110101111010110101111110110110100010011001000010000101010100000111011001001000100101110010101100111000011011101001111101011",
54 => "0100011011100110010010001001101010100001101010001110101001001110100110011011011001000101100011110101000000001011011101111111101011110101010011111111101111101100011110110110011010010110101001010111001001000011011111101111101100010101100111011001001000011100",
55 => "0100110000101010101010000000110010111111001110100010011110110101011011100000001100101100000111011110000100011000011111000000000110100111000100000101001011001100010101100110101110001110111011100100111011101111001010010110110100101000000011111101111000111010",
56 => "1111010100001011011101101010101011100101001010111111011000101110110101010111111010011100011101100111111100000000000110111011111110101011111000011011111001111101100000000000011110011000100111111001011001001101111010001111001001011001101001000110111001010101",
57 => "1001010101000110001001101100100100101010000111110010110110011110001001101000001110110010001010101110000001011000110011011100111010011100011000001011000001110101100010111101000001010010100001110111111011110111100010001110100101011011111000010010100000111000",
58 => "0011000110000001110001000011011111001100110000110100011111100111001000010110010111000110000101011001011001101110100000010100011001011001011111100010101001001100011011111011001110010110001101110001010100001100100111010010000111011100000100101010111000001010",
59 => "1000011101001001100011011000101011110110001011011010001010110111000010101001001001110010110001000001010001010111011001100010010001010001011010011000010000000011011101010111101011101011001010000111101110001101010011000001010110100000100000110011011110011101",
60 => "1111010101101110110110110011011110000110110100011100111111010000111101100101101110111111010001100001101111110111110110000110101000010111111010000110110010010000001011110010111000100111010010100110110010111101011001101011001001111100010000111000001100010011",
61 => "1111110001110001101010001110001000101011111100011111010101110000011000100110000111110100010110100011110100101100001110110011111011001010000100000110000000001010110010100011000011111100001010110111010001100011001010110010000101110011111100001001011111001011",
62 => "1011010100101110000010111110111001010001100000001101010011101000011110110000110100000101101011101000001000101011101111100010101110001000100101000010100110111011011001100111101011110011110010001011010011001010011111110001111010000110010011110101010100111110",
63 => "1100001110000011010101010010010100001110111011110111010001100000101010010111110000110110110111101101001101010000001101110111111010110110001100000011010000000111101110011111000100100110000100001000010010101101010110110101110000111010111001000100100110001111",
64 => "1011110100011000100110110111010110010111011001000000000101010000001100101100001011000110000100111011100000010001110110101010000101001011100101110101101100001001100010010001111111001001011111111001011110010101000100101101101001100100111110110001011001100011",
65 => "1010000111101011110100110010011111101101110100101100000100000000100010110111011111100100000111100111000111101110011010001100011011011010000111110011101110010001011000000110111101111010110001100100000100001110000001000110001000100001110101010001111111110110",
66 => "1100000110110110011111011101110110100011011101000110101010101110001011101110001010111010011100011011100011101011001110101010111010000001011101101111110011000000001001100001111001010101110111001100111101001001101101000011001100110110001110010100000001101111",
67 => "0011000101101000000010110000100011000000101010001000111011110010001001100001111110110011110010010101100000001100000000101000000101001110010001110010111101000000111000011010110110011101000010010101001111100010100110101111000110001010000011101000111001100000",
68 => "0010111111000110111111110101100101010111000001101111000000101110111110111010111001101101110100110110111001100110000101110111011001101111001111101000010011010111111001000101001001010010111100001011000111010010010110000101100111111101111000011111100110100111",
69 => "0100010101110010111100111011011000110101001011010010101001010111100111010001001101110001000000011101011101011110001000011111101111110110100010111100011100101000001000010101011011101110101100110101110001001110010001110011100011110111110111101001111111110111",
70 => "0110100000111011111011000001100111100010010000011101110100100001001010001001101000010100110110011111011110111110110000011000001000011010110010010000100011001011001110100000010000011011111110100011011110110001101000011010011101110111100011010101000110111100",
71 => "0011111111001100110010110010000000011010111011001101110011101111110010001000000101100101101101010111100101110101001111100110101111010110000000011010100100101000111110000001000111111100001000100101110011000111101101100000000101101010111111100110001010010101",
72 => "0110001000101001000001000010111101010000010110000011001111100000011110000011001010011110111000110110001101101100000001010100001001101000001010100010110011000101010101011111101110110011111111111001010010010011101101111110100010101010001101101001100010110010",
73 => "1011110111110001010101110100001000010111110101011001110101011111011000110110001011100101001010010101101011101110111001101001111100000110101001000101100010111100000001001101101001001000011110010100100011000111111000001001101000001000100110011100101011101100",
74 => "1101101011000110001000001010111011010111010001100000111100011110100100100100000100100110011100111111000001110110000110000000101010001100110010100110110001110010001100111110111001101111100111111010111011100001111101110110001111011011110111111100001100110000",
75 => "0000000010010101001100100000001111001100111101011011110000110110101011100111011011100010001010111001011001111011110110101000100001100000111110010011110011100010101101111010111100001110010010111001010111110100111011110101111111100101011111001000001000000000",
76 => "1100101110011101101011001011101111011100101011011101000111100010101110100100011101010110101110110110000100010111000111100010010101010111100001000000100101101111111110110011001001000010010001000010010100001001000010000100010111001011110011010000010000010001",
77 => "1001111110100001101000010010111011001011100000001111111111110000000001110001001000100011000110000100010101001101001110110110000011000011010000111111101001011001110010011100100101110000011100111011001101001101001000011001100010110000100001110000000010011010",
78 => "0110111001001001011011010101110010110000000000010100010100101111110111011000000010001000101011100001100010011000000010011010011101100111010000011100100110101111010110111011010110001011011100001110111110010110010110101110111000110000111011011111111011101111",
79 => "0000000111001110111001100010000001000001010100011100001011111000010001101111100011000011100011101000011000101000110010000110000111000001011100001111110000110010010111101101011101101001010010000101011010011001101111000001001001000110101011010000100101111001",
80 => "0001001100000100110000111101010010010011011110001000100111001111010101010111010011010101111001111100011100100011110011010111010101001010010000010010001110001100101110011110101001000101011001111011101101011111100001110011111000110100001100000001010111011000",
81 => "0001010010001010010110101000011000000010001001101110001101101100101111001011011111111000101011001111100001000100001000101011101011111101011100110110111110011000100010010101010101000000111100100011101011001101000010001101101010111010011001010001100101101010",
82 => "0111110100110001110011001001010110001000000100111100010110010100110101110001110111000010010011011010001000010011010110110111111011110000100010101110110001111100000011101011111010101101110100010011111010101010000101111010100011111010001111000111000001010100",
83 => "1110010111101110100011101100000101001110001111111101001011100111101101101011100001010011010000111101101111110111101001010000111011101111001000111111011000101000001011001010111100111000011111010110010001111110101101000101000100100101111110000010100110100111",
84 => "0011111010100001101001010110110010111011010101100100101001001100111100101101010100111010001110011011011100011000001010000101111010010010100000011101001111000001100011011010111010111000000100100000001101111100010011111000100110100011011101101110010101000111",
85 => "0011100011100010111100100111001101000110001011100000111011000011100111001110010010101110110010001000011101010101111101101000111110110111001100000000000111001000001101110010101110011110011101000101110010001011110011011011101010101001111011101111011001101001",
86 => "0001110011011001011101011001101010010100000011100000011100011010100101001011000011011001110001110011010101010100100110110111011111111011100111010110111111001100001111100110100101011100000010000011000011001010100110111011101111011001000001010111011100101100",
87 => "0101011011100101111010011101001010001000101000101001011101100101001110101001010001100101010100101101000110010011101100100001101100100101010111001001101001011101111100010010001000110011010000000001000010011011000101011000001001110100110000100110010001110101",
88 => "0001010010110101000001011111111000000100000000010101000010111110110000111001000101110011110101000010100111011000010011000011110100110110000100010011000110111101010101100111011100110011111111100101100001100011111000000101101000111100110101111101111110011100",
89 => "1001110011100100010010110110101001110010111001011000010000011100101101110010001011011001100000011111101110001110010100010101000010000100101111100000111100010110111101011001111000011101110000010001001010011100111101011000001001100100110001111110001101110101",
90 => "0010101000010111011001100000000100110010110110010010111001111111110010010101101100000000100111001011111010110101011010010010101011011011010100011011001100100111110010010101110101111011001111010101011010111111001010111001001001100110101011000001100101001001",
91 => "0010111010001010110001000000111001000100011101100010011110100011000010001011111010100000101001111001100001010101110010110001000110010100000010111100111101110010101011011110111001011010011000001010111011000001101111001111101011001111101111100100001000011110",
92 => "1010000110111000110011101010011100001011001100100000001111011010100001001001000110110001000111111011110110100001000100101101110001111010001011100000011110000001110011101011010010101011111101100100010101011100101100011100001011001101111011000011101101011110",
93 => "0011111010000100010010111001111001011111000010111000111111100010001101101100100101101000010110000001001100111011110010100001000101000101000011111100011111111010101000111001110010001100111010001001101001101010101110110000101011010111010101011001010111110100",
94 => "1101011100110100010111101010100101101000000011101000001110000001011000100110010111000001000011100101011110000111100001100000101111000110010100100011100001101001010111001011111110010101001010010100000111101010011111001010111110100111001010000001110110011001",
95 => "1101000011010110110110001101111000000101100110111111001001011101101001100000000010010111101010100010001110100110101000110001101110111111001000011000111100110101111001010010010000100011110101101001001011111001000111100001001101010101010001111100101011101011",
96 => "1100000011110011001111111000001001100111001011111111111101100101010100010111100111100110100110010111101100111100010110111011101110000111001000001110101110010010110001011010110000111011001011000100000000100001000010100100000001101011000101000011011110101100",
97 => "0000111010010000000011110101101011100011111001111010001010110110111101000010100110000101011101101111100111110010000110011000010110111100101111010000011011011011001111010010100000000101110011101101001100111000000101110111000100111000010010010100101100011011",
98 => "0100110111101011110010101101001100001010100101011000101101111001101010010100001101011110000001001101001001111011010111100111010101010010100011110001000000110000101111000011111100001101000101001000100111101111100110000101000101101111110111001110100111000101",
99 => "0011101011010111100110110001100110010101110100110001010110111110110010110010100100101101011110111111011101011000010111111000011111101011001100011101111111000101100101101011011100100001001111000101011011110010110101100010111000101001010100010011001100101011",
100 => "0101000101111111111111111110111100110101010100100111110111001011011111101000010001011001100010010011011010110000011011001010110010011110010001011110001101011110001011101110101110100101000100101010000111111101100101010101110110110110001010000010110110011110"
);

begin

CLOCK_PROGRESS : process
	begin
		Clock<='0';
		wait for clk_period/2;
		Clock<='1';
		wait for clk_period/2;
end process;

tester : process (Clock)
begin

	--test <= ROM_R(0);
	--check <= ROM_C(0);

		if (counter = 100) then
		counter <= 1;
		test <= ROM_R(counter);
		check <= ROM_C(counter);
	else
		counter <= counter + 1;
		test <= ROM_R(counter);
		check <= ROM_C(counter);
	end if;

end process;


checker : process (Clock,result)
begin
	if (result = check) then
		ok <= '1';
	else
		ok <= '0';
	end if;
	
end process;


dut : DecoderBCHE
	port map(
		clock  => Clock,
		input	=> test, --ROM_SINGLEin(0), --test,
		output => result
	);

end architecture;