LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

entity Decoder is
		port(  
		clock  : in std_logic;
		input  : in std_logic_vector(254 downto 0);
		output : out std_logic_vector(254 downto 0)
		);
end entity;

architecture Decoder_arch of Decoder is



type ROM_type is array (1 to 255) of std_logic_vector(7 downto 0);
constant ROM_alpha : ROM_type := ( 1 => "00000001",
2 => "00000010",
3 => "00000100",
4 => "00001000",
5 => "00010000",
6 => "00100000",
7 => "01000000",
8 => "10000000",
9 => "00011101",
10 => "00111010",
11 => "01110100",
12 => "11101000",
13 => "11001101",
14 => "10000111",
15 => "00010011",
16 => "00100110",
17 => "01001100",
18 => "10011000",
19 => "00101101",
20 => "01011010",
21 => "10110100",
22 => "01110101",
23 => "11101010",
24 => "11001001",
25 => "10001111",
26 => "00000011",
27 => "00000110",
28 => "00001100",
29 => "00011000",
30 => "00110000",
31 => "01100000",
32 => "11000000",
33 => "10011101",
34 => "00100111",
35 => "01001110",
36 => "10011100",
37 => "00100101",
38 => "01001010",
39 => "10010100",
40 => "00110101",
41 => "01101010",
42 => "11010100",
43 => "10110101",
44 => "01110111",
45 => "11101110",
46 => "11000001",
47 => "10011111",
48 => "00100011",
49 => "01000110",
50 => "10001100",
51 => "00000101",
52 => "00001010",
53 => "00010100",
54 => "00101000",
55 => "01010000",
56 => "10100000",
57 => "01011101",
58 => "10111010",
59 => "01101001",
60 => "11010010",
61 => "10111001",
62 => "01101111",
63 => "11011110",
64 => "10100001",
65 => "01011111",
66 => "10111110",
67 => "01100001",
68 => "11000010",
69 => "10011001",
70 => "00101111",
71 => "01011110",
72 => "10111100",
73 => "01100101",
74 => "11001010",
75 => "10001001",
76 => "00001111",
77 => "00011110",
78 => "00111100",
79 => "01111000",
80 => "11110000",
81 => "11111101",
82 => "11100111",
83 => "11010011",
84 => "10111011",
85 => "01101011",
86 => "11010110",
87 => "10110001",
88 => "01111111",
89 => "11111110",
90 => "11100001",
91 => "11011111",
92 => "10100011",
93 => "01011011",
94 => "10110110",
95 => "01110001",
96 => "11100010",
97 => "11011001",
98 => "10101111",
99 => "01000011",
100 => "10000110",
101 => "00010001",
102 => "00100010",
103 => "01000100",
104 => "10001000",
105 => "00001101",
106 => "00011010",
107 => "00110100",
108 => "01101000",
109 => "11010000",
110 => "10111101",
111 => "01100111",
112 => "11001110",
113 => "10000001",
114 => "00011111",
115 => "00111110",
116 => "01111100",
117 => "11111000",
118 => "11101101",
119 => "11000111",
120 => "10010011",
121 => "00111011",
122 => "01110110",
123 => "11101100",
124 => "11000101",
125 => "10010111",
126 => "00110011",
127 => "01100110",
128 => "11001100",
129 => "10000101",
130 => "00010111",
131 => "00101110",
132 => "01011100",
133 => "10111000",
134 => "01101101",
135 => "11011010",
136 => "10101001",
137 => "01001111",
138 => "10011110",
139 => "00100001",
140 => "01000010",
141 => "10000100",
142 => "00010101",
143 => "00101010",
144 => "01010100",
145 => "10101000",
146 => "01001101",
147 => "10011010",
148 => "00101001",
149 => "01010010",
150 => "10100100",
151 => "01010101",
152 => "10101010",
153 => "01001001",
154 => "10010010",
155 => "00111001",
156 => "01110010",
157 => "11100100",
158 => "11010101",
159 => "10110111",
160 => "01110011",
161 => "11100110",
162 => "11010001",
163 => "10111111",
164 => "01100011",
165 => "11000110",
166 => "10010001",
167 => "00111111",
168 => "01111110",
169 => "11111100",
170 => "11100101",
171 => "11010111",
172 => "10110011",
173 => "01111011",
174 => "11110110",
175 => "11110001",
176 => "11111111",
177 => "11100011",
178 => "11011011",
179 => "10101011",
180 => "01001011",
181 => "10010110",
182 => "00110001",
183 => "01100010",
184 => "11000100",
185 => "10010101",
186 => "00110111",
187 => "01101110",
188 => "11011100",
189 => "10100101",
190 => "01010111",
191 => "10101110",
192 => "01000001",
193 => "10000010",
194 => "00011001",
195 => "00110010",
196 => "01100100",
197 => "11001000",
198 => "10001101",
199 => "00000111",
200 => "00001110",
201 => "00011100",
202 => "00111000",
203 => "01110000",
204 => "11100000",
205 => "11011101",
206 => "10100111",
207 => "01010011",
208 => "10100110",
209 => "01010001",
210 => "10100010",
211 => "01011001",
212 => "10110010",
213 => "01111001",
214 => "11110010",
215 => "11111001",
216 => "11101111",
217 => "11000011",
218 => "10011011",
219 => "00101011",
220 => "01010110",
221 => "10101100",
222 => "01000101",
223 => "10001010",
224 => "00001001",
225 => "00010010",
226 => "00100100",
227 => "01001000",
228 => "10010000",
229 => "00111101",
230 => "01111010",
231 => "11110100",
232 => "11110101",
233 => "11110111",
234 => "11110011",
235 => "11111011",
236 => "11101011",
237 => "11001011",
238 => "10001011",
239 => "00001011",
240 => "00010110",
241 => "00101100",
242 => "01011000",
243 => "10110000",
244 => "01111101",
245 => "11111010",
246 => "11101001",
247 => "11001111",
248 => "10000011",
249 => "00011011",
250 => "00110110",
251 => "01101100",
252 => "11011000",
253 => "10101101",
254 => "01000111",
255 => "10001110");

type ROM_type2 is array (1 to 255) of integer;
constant ROM_alphaInv : ROM_type2 := ( 1 => 0,
2 => 1,
3 => 25,
4 => 2,
5 => 50,
6 => 26,
7 => 198,
8 => 3,
9 => 223,
10 => 51,
11 => 238,
12 => 27,
13 => 104,
14 => 199,
15 => 75,
16 => 4,
17 => 100,
18 => 224,
19 => 14,
20 => 52,
21 => 141,
22 => 239,
23 => 129,
24 => 28,
25 => 193,
26 => 105,
27 => 248,
28 => 200,
29 => 8,
30 => 76,
31 => 113,
32 => 5,
33 => 138,
34 => 101,
35 => 47,
36 => 225,
37 => 36,
38 => 15,
39 => 33,
40 => 53,
41 => 147,
42 => 142,
43 => 218,
44 => 240,
45 => 18,
46 => 130,
47 => 69,
48 => 29,
49 => 181,
50 => 194,
51 => 125,
52 => 106,
53 => 39,
54 => 249,
55 => 185,
56 => 201,
57 => 154,
58 => 9,
59 => 120,
60 => 77,
61 => 228,
62 => 114,
63 => 166,
64 => 6,
65 => 191,
66 => 139,
67 => 98,
68 => 102,
69 => 221,
70 => 48,
71 => 253,
72 => 226,
73 => 152,
74 => 37,
75 => 179,
76 => 16,
77 => 145,
78 => 34,
79 => 136,
80 => 54,
81 => 208,
82 => 148,
83 => 206,
84 => 143,
85 => 150,
86 => 219,
87 => 189,
88 => 241,
89 => 210,
90 => 19,
91 => 92,
92 => 131,
93 => 56,
94 => 70,
95 => 64,
96 => 30,
97 => 66,
98 => 182,
99 => 163,
100 => 195,
101 => 72,
102 => 126,
103 => 110,
104 => 107,
105 => 58,
106 => 40,
107 => 84,
108 => 250,
109 => 133,
110 => 186,
111 => 61,
112 => 202,
113 => 94,
114 => 155,
115 => 159,
116 => 10,
117 => 21,
118 => 121,
119 => 43,
120 => 78,
121 => 212,
122 => 229,
123 => 172,
124 => 115,
125 => 243,
126 => 167,
127 => 87,
128 => 7,
129 => 112,
130 => 192,
131 => 247,
132 => 140,
133 => 128,
134 => 99,
135 => 13,
136 => 103,
137 => 74,
138 => 222,
139 => 237,
140 => 49,
141 => 197,
142 => 254,
143 => 24,
144 => 227,
145 => 165,
146 => 153,
147 => 119,
148 => 38,
149 => 184,
150 => 180,
151 => 124,
152 => 17,
153 => 68,
154 => 146,
155 => 217,
156 => 35,
157 => 32,
158 => 137,
159 => 46,
160 => 55,
161 => 63,
162 => 209,
163 => 91,
164 => 149,
165 => 188,
166 => 207,
167 => 205,
168 => 144,
169 => 135,
170 => 151,
171 => 178,
172 => 220,
173 => 252,
174 => 190,
175 => 97,
176 => 242,
177 => 86,
178 => 211,
179 => 171,
180 => 20,
181 => 42,
182 => 93,
183 => 158,
184 => 132,
185 => 60,
186 => 57,
187 => 83,
188 => 71,
189 => 109,
190 => 65,
191 => 162,
192 => 31,
193 => 45,
194 => 67,
195 => 216,
196 => 183,
197 => 123,
198 => 164,
199 => 118,
200 => 196,
201 => 23,
202 => 73,
203 => 236,
204 => 127,
205 => 12,
206 => 111,
207 => 246,
208 => 108,
209 => 161,
210 => 59,
211 => 82,
212 => 41,
213 => 157,
214 => 85,
215 => 170,
216 => 251,
217 => 96,
218 => 134,
219 => 177,
220 => 187,
221 => 204,
222 => 62,
223 => 90,
224 => 203,
225 => 89,
226 => 95,
227 => 176,
228 => 156,
229 => 169,
230 => 160,
231 => 81,
232 => 11,
233 => 245,
234 => 22,
235 => 235,
236 => 122,
237 => 117,
238 => 44,
239 => 215,
240 => 79,
241 => 174,
242 => 213,
243 => 233,
244 => 230,
245 => 231,
246 => 173,
247 => 232,
248 => 116,
249 => 214,
250 => 244,
251 => 234,
252 => 168,
253 => 80,
254 => 88,
255 => 175);





type ROM_type3 is array (0 to 254) of integer;
constant ROM_yFirstMatch : ROM_type3 := ( 0 => 85,
1 => 11,
2 => 22,
3 => 18,
4 => 44,
5 => 0,
6 => 36,
7 => 54,
8 => 88,
9 => 0,
10 => 0,
11 => 0,
12 => 72,
13 => 128,
14 => 108,
15 => 0,
16 => 95,
17 => 119,
18 => 0,
19 => 75,
20 => 0,
21 => 0,
22 => 0,
23 => 24,
24 => 135,
25 => 114,
26 => 1,
27 => 118,
28 => 67,
29 => 0,
30 => 0,
31 => 10,
32 => 97,
33 => 0,
34 => 51,
35 => 78,
36 => 0,
37 => 89,
38 => 143,
39 => 0,
40 => 0,
41 => 94,
42 => 0,
43 => 0,
44 => 0,
45 => 91,
46 => 48,
47 => 0,
48 => 15,
49 => 124,
50 => 77,
51 => 123,
52 => 2,
53 => 0,
54 => 73,
55 => 0,
56 => 134,
57 => 0,
58 => 0,
59 => 155,
60 => 0,
61 => 0,
62 => 20,
63 => 0,
64 => 125,
65 => 0,
66 => 0,
67 => 32,
68 => 102,
69 => 0,
70 => 156,
71 => 0,
72 => 0,
73 => 86,
74 => 151,
75 => 116,
76 => 31,
77 => 0,
78 => 0,
79 => 0,
80 => 0,
81 => 0,
82 => 149,
83 => 0,
84 => 0,
85 => 17,
86 => 0,
87 => 0,
88 => 0,
89 => 0,
90 => 163,
91 => 0,
92 => 96,
93 => 0,
94 => 0,
95 => 0,
96 => 30,
97 => 0,
98 => 105,
99 => 148,
100 => 154,
101 => 0,
102 => 111,
103 => 115,
104 => 4,
105 => 142,
106 => 0,
107 => 0,
108 => 146,
109 => 0,
110 => 0,
111 => 19,
112 => 13,
113 => 129,
114 => 0,
115 => 0,
116 => 0,
117 => 0,
118 => 55,
119 => 7,
120 => 0,
121 => 0,
122 => 0,
123 => 152,
124 => 40,
125 => 0,
126 => 0,
127 => 171,
128 => 133,
129 => 9,
130 => 0,
131 => 27,
132 => 0,
133 => 0,
134 => 64,
135 => 0,
136 => 187,
137 => 165,
138 => 0,
139 => 12,
140 => 57,
141 => 59,
142 => 0,
143 => 5,
144 => 0,
145 => 39,
146 => 172,
147 => 0,
148 => 47,
149 => 0,
150 => 173,
151 => 0,
152 => 62,
153 => 189,
154 => 0,
155 => 0,
156 => 0,
157 => 205,
158 => 0,
159 => 0,
160 => 0,
161 => 16,
162 => 0,
163 => 0,
164 => 43,
165 => 58,
166 => 0,
167 => 0,
168 => 0,
169 => 0,
170 => 34,
171 => 0,
172 => 0,
173 => 0,
174 => 0,
175 => 0,
176 => 0,
177 => 74,
178 => 0,
179 => 185,
180 => 71,
181 => 0,
182 => 0,
183 => 46,
184 => 192,
185 => 0,
186 => 0,
187 => 56,
188 => 0,
189 => 76,
190 => 0,
191 => 213,
192 => 60,
193 => 52,
194 => 0,
195 => 0,
196 => 210,
197 => 6,
198 => 41,
199 => 69,
200 => 53,
201 => 0,
202 => 0,
203 => 0,
204 => 222,
205 => 0,
206 => 230,
207 => 0,
208 => 8,
209 => 0,
210 => 29,
211 => 0,
212 => 0,
213 => 0,
214 => 0,
215 => 0,
216 => 37,
217 => 220,
218 => 0,
219 => 23,
220 => 0,
221 => 28,
222 => 38,
223 => 234,
224 => 26,
225 => 0,
226 => 3,
227 => 65,
228 => 0,
229 => 0,
230 => 0,
231 => 0,
232 => 0,
233 => 0,
234 => 0,
235 => 0,
236 => 110,
237 => 98,
238 => 14,
239 => 117,
240 => 0,
241 => 81,
242 => 0,
243 => 0,
244 => 0,
245 => 0,
246 => 49,
247 => 61,
248 => 80,
249 => 0,
250 => 0,
251 => 93,
252 => 0,
253 => 79,
254 => 87
);


constant ROM_ySecondMatch : ROM_type3 := ( 0 => 170,
1 => 245,
2 => 235,
3 => 240,
4 => 215,
5 => 0,
6 => 225,
7 => 208,
8 => 175,
9 => 0,
10 => 0,
11 => 0,
12 => 195,
13 => 140,
14 => 161,
15 => 0,
16 => 176,
17 => 153,
18 => 0,
19 => 199,
20 => 0,
21 => 0,
22 => 0,
23 => 254,
24 => 144,
25 => 166,
26 => 25,
27 => 164,
28 => 216,
29 => 0,
30 => 0,
31 => 21,
32 => 190,
33 => 0,
34 => 238,
35 => 212,
36 => 0,
37 => 203,
38 => 150,
39 => 0,
40 => 0,
41 => 202,
42 => 0,
43 => 0,
44 => 0,
45 => 209,
46 => 253,
47 => 0,
48 => 33,
49 => 180,
50 => 228,
51 => 183,
52 => 50,
53 => 0,
54 => 236,
55 => 0,
56 => 177,
57 => 0,
58 => 0,
59 => 159,
60 => 0,
61 => 0,
62 => 42,
63 => 0,
64 => 194,
65 => 0,
66 => 0,
67 => 35,
68 => 221,
69 => 0,
70 => 169,
71 => 0,
72 => 0,
73 => 242,
74 => 178,
75 => 214,
76 => 45,
77 => 0,
78 => 0,
79 => 0,
80 => 0,
81 => 0,
82 => 188,
83 => 0,
84 => 0,
85 => 68,
86 => 0,
87 => 0,
88 => 0,
89 => 0,
90 => 182,
91 => 0,
92 => 251,
93 => 0,
94 => 0,
95 => 0,
96 => 66,
97 => 0,
98 => 248,
99 => 206,
100 => 201,
101 => 0,
102 => 246,
103 => 243,
104 => 100,
105 => 218,
106 => 0,
107 => 0,
108 => 217,
109 => 0,
110 => 0,
111 => 92,
112 => 99,
113 => 239,
114 => 0,
115 => 0,
116 => 0,
117 => 0,
118 => 63,
119 => 112,
120 => 0,
121 => 0,
122 => 0,
123 => 226,
124 => 84,
125 => 0,
126 => 0,
127 => 211,
128 => 250,
129 => 120,
130 => 0,
131 => 104,
132 => 0,
133 => 0,
134 => 70,
135 => 0,
136 => 204,
137 => 227,
138 => 0,
139 => 127,
140 => 83,
141 => 82,
142 => 0,
143 => 138,
144 => 0,
145 => 106,
146 => 229,
147 => 0,
148 => 101,
149 => 0,
150 => 232,
151 => 0,
152 => 90,
153 => 219,
154 => 0,
155 => 0,
156 => 0,
157 => 207,
158 => 0,
159 => 0,
160 => 0,
161 => 145,
162 => 0,
163 => 0,
164 => 121,
165 => 107,
166 => 0,
167 => 0,
168 => 0,
169 => 0,
170 => 136,
171 => 0,
172 => 0,
173 => 0,
174 => 0,
175 => 0,
176 => 0,
177 => 103,
178 => 0,
179 => 249,
180 => 109,
181 => 0,
182 => 0,
183 => 137,
184 => 247,
185 => 0,
186 => 0,
187 => 131,
188 => 0,
189 => 113,
190 => 0,
191 => 233,
192 => 132,
193 => 141,
194 => 0,
195 => 0,
196 => 241,
197 => 191,
198 => 157,
199 => 130,
200 => 147,
201 => 0,
202 => 0,
203 => 0,
204 => 237,
205 => 0,
206 => 231,
207 => 0,
208 => 200,
209 => 0,
210 => 181,
211 => 0,
212 => 0,
213 => 0,
214 => 0,
215 => 0,
216 => 179,
217 => 252,
218 => 0,
219 => 196,
220 => 0,
221 => 193,
222 => 184,
223 => 244,
224 => 198,
225 => 0,
226 => 223,
227 => 162,
228 => 0,
229 => 0,
230 => 0,
231 => 0,
232 => 0,
233 => 0,
234 => 0,
235 => 0,
236 => 126,
237 => 139,
238 => 224,
239 => 122,
240 => 0,
241 => 160,
242 => 0,
243 => 0,
244 => 0,
245 => 0,
246 => 197,
247 => 186,
248 => 168,
249 => 0,
250 => 0,
251 => 158,
252 => 0,
253 => 174,
254 => 167
);

type ROM_type4 is array (0 to 255) of std_logic_vector(254 downto 0);
constant ROM_E : ROM_type4 := ( 
0 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
1 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001",
2 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010",
3 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100",
4 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000",
5 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000",
6 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000",
7 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000",
8 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000",
9 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000",
10 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000",
11 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000",
12 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000",
13 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000",
14 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000",
15 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000",
16 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000",
17 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000",
18 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000",
19 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000",
20 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000",
21 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000",
22 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000",
23 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000",
24 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000",
25 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000",
26 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000",
27 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000",
28 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000",
29 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000",
30 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000",
31 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000",
32 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000",
33 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000",
34 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000",
35 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000",
36 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000",
37 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000",
38 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000",
39 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000",
40 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000",
41 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000",
42 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000",
43 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000",
44 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000",
45 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000",
46 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000",
47 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000",
48 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000",
49 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000",
50 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000",
51 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000",
52 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000",
53 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000",
54 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000",
55 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000",
56 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000",
57 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000",
58 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000",
59 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000",
60 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000",
61 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000",
62 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000",
63 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000",
64 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000",
65 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000",
66 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000",
67 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000",
68 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000",
69 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000",
70 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000",
71 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000",
72 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000",
73 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000",
74 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000",
75 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000",
76 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000",
77 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000",
78 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000",
79 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000",
80 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000",
81 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000",
82 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000",
83 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000",
84 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000",
85 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
86 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
87 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
88 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
89 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
90 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
91 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
92 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
93 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
94 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
95 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
96 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
97 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
98 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
99 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
100 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
101 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
102 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
103 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
104 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
105 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
106 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
107 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
108 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
109 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
110 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
111 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
112 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
113 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
114 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
115 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
116 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
117 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
118 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
119 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
120 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
121 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
122 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
123 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
124 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
125 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
126 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
127 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
128 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
129 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
130 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
131 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
132 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
133 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
134 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
135 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
136 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
137 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
138 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
139 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
140 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
141 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
142 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
143 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
144 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
145 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
146 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
147 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
148 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
149 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
150 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
151 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
152 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
153 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
154 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
155 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
156 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
157 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
158 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
159 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
160 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
161 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
162 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
163 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
164 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
165 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
166 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
167 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
168 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
169 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
170 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
171 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
172 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
173 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
174 => "000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
175 => "000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
176 => "000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
177 => "000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
178 => "000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
179 => "000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
180 => "000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
181 => "000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
182 => "000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
183 => "000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
184 => "000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
185 => "000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
186 => "000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
187 => "000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
188 => "000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
189 => "000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
190 => "000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
191 => "000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
192 => "000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
193 => "000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
194 => "000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
195 => "000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
196 => "000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
197 => "000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
198 => "000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
199 => "000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
200 => "000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
201 => "000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
202 => "000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
203 => "000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
204 => "000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
205 => "000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
206 => "000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
207 => "000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
208 => "000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
209 => "000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
210 => "000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
211 => "000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
212 => "000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
213 => "000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
214 => "000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
215 => "000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
216 => "000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
217 => "000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
218 => "000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
219 => "000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
220 => "000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
221 => "000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
222 => "000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
223 => "000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
224 => "000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
225 => "000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
226 => "000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
227 => "000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
228 => "000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
229 => "000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
230 => "000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
231 => "000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
232 => "000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
233 => "000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
234 => "000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
235 => "000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
236 => "000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
237 => "000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
238 => "000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
239 => "000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
240 => "000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
241 => "000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
242 => "000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
243 => "000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
244 => "000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
245 => "000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
246 => "000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
247 => "000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
248 => "000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
249 => "000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
250 => "000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
251 => "000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
252 => "000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
253 => "001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
254 => "010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000",
255 => "100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000"
);


type ROM_type5 is array (-765 to 765) of integer;
constant ROM_MOD : ROM_type5 := ( -765 => 0,
-764 => 1,
-763 => 2,
-762 => 3,
-761 => 4,
-760 => 5,
-759 => 6,
-758 => 7,
-757 => 8,
-756 => 9,
-755 => 10,
-754 => 11,
-753 => 12,
-752 => 13,
-751 => 14,
-750 => 15,
-749 => 16,
-748 => 17,
-747 => 18,
-746 => 19,
-745 => 20,
-744 => 21,
-743 => 22,
-742 => 23,
-741 => 24,
-740 => 25,
-739 => 26,
-738 => 27,
-737 => 28,
-736 => 29,
-735 => 30,
-734 => 31,
-733 => 32,
-732 => 33,
-731 => 34,
-730 => 35,
-729 => 36,
-728 => 37,
-727 => 38,
-726 => 39,
-725 => 40,
-724 => 41,
-723 => 42,
-722 => 43,
-721 => 44,
-720 => 45,
-719 => 46,
-718 => 47,
-717 => 48,
-716 => 49,
-715 => 50,
-714 => 51,
-713 => 52,
-712 => 53,
-711 => 54,
-710 => 55,
-709 => 56,
-708 => 57,
-707 => 58,
-706 => 59,
-705 => 60,
-704 => 61,
-703 => 62,
-702 => 63,
-701 => 64,
-700 => 65,
-699 => 66,
-698 => 67,
-697 => 68,
-696 => 69,
-695 => 70,
-694 => 71,
-693 => 72,
-692 => 73,
-691 => 74,
-690 => 75,
-689 => 76,
-688 => 77,
-687 => 78,
-686 => 79,
-685 => 80,
-684 => 81,
-683 => 82,
-682 => 83,
-681 => 84,
-680 => 85,
-679 => 86,
-678 => 87,
-677 => 88,
-676 => 89,
-675 => 90,
-674 => 91,
-673 => 92,
-672 => 93,
-671 => 94,
-670 => 95,
-669 => 96,
-668 => 97,
-667 => 98,
-666 => 99,
-665 => 100,
-664 => 101,
-663 => 102,
-662 => 103,
-661 => 104,
-660 => 105,
-659 => 106,
-658 => 107,
-657 => 108,
-656 => 109,
-655 => 110,
-654 => 111,
-653 => 112,
-652 => 113,
-651 => 114,
-650 => 115,
-649 => 116,
-648 => 117,
-647 => 118,
-646 => 119,
-645 => 120,
-644 => 121,
-643 => 122,
-642 => 123,
-641 => 124,
-640 => 125,
-639 => 126,
-638 => 127,
-637 => 128,
-636 => 129,
-635 => 130,
-634 => 131,
-633 => 132,
-632 => 133,
-631 => 134,
-630 => 135,
-629 => 136,
-628 => 137,
-627 => 138,
-626 => 139,
-625 => 140,
-624 => 141,
-623 => 142,
-622 => 143,
-621 => 144,
-620 => 145,
-619 => 146,
-618 => 147,
-617 => 148,
-616 => 149,
-615 => 150,
-614 => 151,
-613 => 152,
-612 => 153,
-611 => 154,
-610 => 155,
-609 => 156,
-608 => 157,
-607 => 158,
-606 => 159,
-605 => 160,
-604 => 161,
-603 => 162,
-602 => 163,
-601 => 164,
-600 => 165,
-599 => 166,
-598 => 167,
-597 => 168,
-596 => 169,
-595 => 170,
-594 => 171,
-593 => 172,
-592 => 173,
-591 => 174,
-590 => 175,
-589 => 176,
-588 => 177,
-587 => 178,
-586 => 179,
-585 => 180,
-584 => 181,
-583 => 182,
-582 => 183,
-581 => 184,
-580 => 185,
-579 => 186,
-578 => 187,
-577 => 188,
-576 => 189,
-575 => 190,
-574 => 191,
-573 => 192,
-572 => 193,
-571 => 194,
-570 => 195,
-569 => 196,
-568 => 197,
-567 => 198,
-566 => 199,
-565 => 200,
-564 => 201,
-563 => 202,
-562 => 203,
-561 => 204,
-560 => 205,
-559 => 206,
-558 => 207,
-557 => 208,
-556 => 209,
-555 => 210,
-554 => 211,
-553 => 212,
-552 => 213,
-551 => 214,
-550 => 215,
-549 => 216,
-548 => 217,
-547 => 218,
-546 => 219,
-545 => 220,
-544 => 221,
-543 => 222,
-542 => 223,
-541 => 224,
-540 => 225,
-539 => 226,
-538 => 227,
-537 => 228,
-536 => 229,
-535 => 230,
-534 => 231,
-533 => 232,
-532 => 233,
-531 => 234,
-530 => 235,
-529 => 236,
-528 => 237,
-527 => 238,
-526 => 239,
-525 => 240,
-524 => 241,
-523 => 242,
-522 => 243,
-521 => 244,
-520 => 245,
-519 => 246,
-518 => 247,
-517 => 248,
-516 => 249,
-515 => 250,
-514 => 251,
-513 => 252,
-512 => 253,
-511 => 254,
-510 => 0,
-509 => 1,
-508 => 2,
-507 => 3,
-506 => 4,
-505 => 5,
-504 => 6,
-503 => 7,
-502 => 8,
-501 => 9,
-500 => 10,
-499 => 11,
-498 => 12,
-497 => 13,
-496 => 14,
-495 => 15,
-494 => 16,
-493 => 17,
-492 => 18,
-491 => 19,
-490 => 20,
-489 => 21,
-488 => 22,
-487 => 23,
-486 => 24,
-485 => 25,
-484 => 26,
-483 => 27,
-482 => 28,
-481 => 29,
-480 => 30,
-479 => 31,
-478 => 32,
-477 => 33,
-476 => 34,
-475 => 35,
-474 => 36,
-473 => 37,
-472 => 38,
-471 => 39,
-470 => 40,
-469 => 41,
-468 => 42,
-467 => 43,
-466 => 44,
-465 => 45,
-464 => 46,
-463 => 47,
-462 => 48,
-461 => 49,
-460 => 50,
-459 => 51,
-458 => 52,
-457 => 53,
-456 => 54,
-455 => 55,
-454 => 56,
-453 => 57,
-452 => 58,
-451 => 59,
-450 => 60,
-449 => 61,
-448 => 62,
-447 => 63,
-446 => 64,
-445 => 65,
-444 => 66,
-443 => 67,
-442 => 68,
-441 => 69,
-440 => 70,
-439 => 71,
-438 => 72,
-437 => 73,
-436 => 74,
-435 => 75,
-434 => 76,
-433 => 77,
-432 => 78,
-431 => 79,
-430 => 80,
-429 => 81,
-428 => 82,
-427 => 83,
-426 => 84,
-425 => 85,
-424 => 86,
-423 => 87,
-422 => 88,
-421 => 89,
-420 => 90,
-419 => 91,
-418 => 92,
-417 => 93,
-416 => 94,
-415 => 95,
-414 => 96,
-413 => 97,
-412 => 98,
-411 => 99,
-410 => 100,
-409 => 101,
-408 => 102,
-407 => 103,
-406 => 104,
-405 => 105,
-404 => 106,
-403 => 107,
-402 => 108,
-401 => 109,
-400 => 110,
-399 => 111,
-398 => 112,
-397 => 113,
-396 => 114,
-395 => 115,
-394 => 116,
-393 => 117,
-392 => 118,
-391 => 119,
-390 => 120,
-389 => 121,
-388 => 122,
-387 => 123,
-386 => 124,
-385 => 125,
-384 => 126,
-383 => 127,
-382 => 128,
-381 => 129,
-380 => 130,
-379 => 131,
-378 => 132,
-377 => 133,
-376 => 134,
-375 => 135,
-374 => 136,
-373 => 137,
-372 => 138,
-371 => 139,
-370 => 140,
-369 => 141,
-368 => 142,
-367 => 143,
-366 => 144,
-365 => 145,
-364 => 146,
-363 => 147,
-362 => 148,
-361 => 149,
-360 => 150,
-359 => 151,
-358 => 152,
-357 => 153,
-356 => 154,
-355 => 155,
-354 => 156,
-353 => 157,
-352 => 158,
-351 => 159,
-350 => 160,
-349 => 161,
-348 => 162,
-347 => 163,
-346 => 164,
-345 => 165,
-344 => 166,
-343 => 167,
-342 => 168,
-341 => 169,
-340 => 170,
-339 => 171,
-338 => 172,
-337 => 173,
-336 => 174,
-335 => 175,
-334 => 176,
-333 => 177,
-332 => 178,
-331 => 179,
-330 => 180,
-329 => 181,
-328 => 182,
-327 => 183,
-326 => 184,
-325 => 185,
-324 => 186,
-323 => 187,
-322 => 188,
-321 => 189,
-320 => 190,
-319 => 191,
-318 => 192,
-317 => 193,
-316 => 194,
-315 => 195,
-314 => 196,
-313 => 197,
-312 => 198,
-311 => 199,
-310 => 200,
-309 => 201,
-308 => 202,
-307 => 203,
-306 => 204,
-305 => 205,
-304 => 206,
-303 => 207,
-302 => 208,
-301 => 209,
-300 => 210,
-299 => 211,
-298 => 212,
-297 => 213,
-296 => 214,
-295 => 215,
-294 => 216,
-293 => 217,
-292 => 218,
-291 => 219,
-290 => 220,
-289 => 221,
-288 => 222,
-287 => 223,
-286 => 224,
-285 => 225,
-284 => 226,
-283 => 227,
-282 => 228,
-281 => 229,
-280 => 230,
-279 => 231,
-278 => 232,
-277 => 233,
-276 => 234,
-275 => 235,
-274 => 236,
-273 => 237,
-272 => 238,
-271 => 239,
-270 => 240,
-269 => 241,
-268 => 242,
-267 => 243,
-266 => 244,
-265 => 245,
-264 => 246,
-263 => 247,
-262 => 248,
-261 => 249,
-260 => 250,
-259 => 251,
-258 => 252,
-257 => 253,
-256 => 254,
-255 => 0,
-254 => 1,
-253 => 2,
-252 => 3,
-251 => 4,
-250 => 5,
-249 => 6,
-248 => 7,
-247 => 8,
-246 => 9,
-245 => 10,
-244 => 11,
-243 => 12,
-242 => 13,
-241 => 14,
-240 => 15,
-239 => 16,
-238 => 17,
-237 => 18,
-236 => 19,
-235 => 20,
-234 => 21,
-233 => 22,
-232 => 23,
-231 => 24,
-230 => 25,
-229 => 26,
-228 => 27,
-227 => 28,
-226 => 29,
-225 => 30,
-224 => 31,
-223 => 32,
-222 => 33,
-221 => 34,
-220 => 35,
-219 => 36,
-218 => 37,
-217 => 38,
-216 => 39,
-215 => 40,
-214 => 41,
-213 => 42,
-212 => 43,
-211 => 44,
-210 => 45,
-209 => 46,
-208 => 47,
-207 => 48,
-206 => 49,
-205 => 50,
-204 => 51,
-203 => 52,
-202 => 53,
-201 => 54,
-200 => 55,
-199 => 56,
-198 => 57,
-197 => 58,
-196 => 59,
-195 => 60,
-194 => 61,
-193 => 62,
-192 => 63,
-191 => 64,
-190 => 65,
-189 => 66,
-188 => 67,
-187 => 68,
-186 => 69,
-185 => 70,
-184 => 71,
-183 => 72,
-182 => 73,
-181 => 74,
-180 => 75,
-179 => 76,
-178 => 77,
-177 => 78,
-176 => 79,
-175 => 80,
-174 => 81,
-173 => 82,
-172 => 83,
-171 => 84,
-170 => 85,
-169 => 86,
-168 => 87,
-167 => 88,
-166 => 89,
-165 => 90,
-164 => 91,
-163 => 92,
-162 => 93,
-161 => 94,
-160 => 95,
-159 => 96,
-158 => 97,
-157 => 98,
-156 => 99,
-155 => 100,
-154 => 101,
-153 => 102,
-152 => 103,
-151 => 104,
-150 => 105,
-149 => 106,
-148 => 107,
-147 => 108,
-146 => 109,
-145 => 110,
-144 => 111,
-143 => 112,
-142 => 113,
-141 => 114,
-140 => 115,
-139 => 116,
-138 => 117,
-137 => 118,
-136 => 119,
-135 => 120,
-134 => 121,
-133 => 122,
-132 => 123,
-131 => 124,
-130 => 125,
-129 => 126,
-128 => 127,
-127 => 128,
-126 => 129,
-125 => 130,
-124 => 131,
-123 => 132,
-122 => 133,
-121 => 134,
-120 => 135,
-119 => 136,
-118 => 137,
-117 => 138,
-116 => 139,
-115 => 140,
-114 => 141,
-113 => 142,
-112 => 143,
-111 => 144,
-110 => 145,
-109 => 146,
-108 => 147,
-107 => 148,
-106 => 149,
-105 => 150,
-104 => 151,
-103 => 152,
-102 => 153,
-101 => 154,
-100 => 155,
-99 => 156,
-98 => 157,
-97 => 158,
-96 => 159,
-95 => 160,
-94 => 161,
-93 => 162,
-92 => 163,
-91 => 164,
-90 => 165,
-89 => 166,
-88 => 167,
-87 => 168,
-86 => 169,
-85 => 170,
-84 => 171,
-83 => 172,
-82 => 173,
-81 => 174,
-80 => 175,
-79 => 176,
-78 => 177,
-77 => 178,
-76 => 179,
-75 => 180,
-74 => 181,
-73 => 182,
-72 => 183,
-71 => 184,
-70 => 185,
-69 => 186,
-68 => 187,
-67 => 188,
-66 => 189,
-65 => 190,
-64 => 191,
-63 => 192,
-62 => 193,
-61 => 194,
-60 => 195,
-59 => 196,
-58 => 197,
-57 => 198,
-56 => 199,
-55 => 200,
-54 => 201,
-53 => 202,
-52 => 203,
-51 => 204,
-50 => 205,
-49 => 206,
-48 => 207,
-47 => 208,
-46 => 209,
-45 => 210,
-44 => 211,
-43 => 212,
-42 => 213,
-41 => 214,
-40 => 215,
-39 => 216,
-38 => 217,
-37 => 218,
-36 => 219,
-35 => 220,
-34 => 221,
-33 => 222,
-32 => 223,
-31 => 224,
-30 => 225,
-29 => 226,
-28 => 227,
-27 => 228,
-26 => 229,
-25 => 230,
-24 => 231,
-23 => 232,
-22 => 233,
-21 => 234,
-20 => 235,
-19 => 236,
-18 => 237,
-17 => 238,
-16 => 239,
-15 => 240,
-14 => 241,
-13 => 242,
-12 => 243,
-11 => 244,
-10 => 245,
-9 => 246,
-8 => 247,
-7 => 248,
-6 => 249,
-5 => 250,
-4 => 251,
-3 => 252,
-2 => 253,
-1 => 254,
0 => 0,
1 => 1,
2 => 2,
3 => 3,
4 => 4,
5 => 5,
6 => 6,
7 => 7,
8 => 8,
9 => 9,
10 => 10,
11 => 11,
12 => 12,
13 => 13,
14 => 14,
15 => 15,
16 => 16,
17 => 17,
18 => 18,
19 => 19,
20 => 20,
21 => 21,
22 => 22,
23 => 23,
24 => 24,
25 => 25,
26 => 26,
27 => 27,
28 => 28,
29 => 29,
30 => 30,
31 => 31,
32 => 32,
33 => 33,
34 => 34,
35 => 35,
36 => 36,
37 => 37,
38 => 38,
39 => 39,
40 => 40,
41 => 41,
42 => 42,
43 => 43,
44 => 44,
45 => 45,
46 => 46,
47 => 47,
48 => 48,
49 => 49,
50 => 50,
51 => 51,
52 => 52,
53 => 53,
54 => 54,
55 => 55,
56 => 56,
57 => 57,
58 => 58,
59 => 59,
60 => 60,
61 => 61,
62 => 62,
63 => 63,
64 => 64,
65 => 65,
66 => 66,
67 => 67,
68 => 68,
69 => 69,
70 => 70,
71 => 71,
72 => 72,
73 => 73,
74 => 74,
75 => 75,
76 => 76,
77 => 77,
78 => 78,
79 => 79,
80 => 80,
81 => 81,
82 => 82,
83 => 83,
84 => 84,
85 => 85,
86 => 86,
87 => 87,
88 => 88,
89 => 89,
90 => 90,
91 => 91,
92 => 92,
93 => 93,
94 => 94,
95 => 95,
96 => 96,
97 => 97,
98 => 98,
99 => 99,
100 => 100,
101 => 101,
102 => 102,
103 => 103,
104 => 104,
105 => 105,
106 => 106,
107 => 107,
108 => 108,
109 => 109,
110 => 110,
111 => 111,
112 => 112,
113 => 113,
114 => 114,
115 => 115,
116 => 116,
117 => 117,
118 => 118,
119 => 119,
120 => 120,
121 => 121,
122 => 122,
123 => 123,
124 => 124,
125 => 125,
126 => 126,
127 => 127,
128 => 128,
129 => 129,
130 => 130,
131 => 131,
132 => 132,
133 => 133,
134 => 134,
135 => 135,
136 => 136,
137 => 137,
138 => 138,
139 => 139,
140 => 140,
141 => 141,
142 => 142,
143 => 143,
144 => 144,
145 => 145,
146 => 146,
147 => 147,
148 => 148,
149 => 149,
150 => 150,
151 => 151,
152 => 152,
153 => 153,
154 => 154,
155 => 155,
156 => 156,
157 => 157,
158 => 158,
159 => 159,
160 => 160,
161 => 161,
162 => 162,
163 => 163,
164 => 164,
165 => 165,
166 => 166,
167 => 167,
168 => 168,
169 => 169,
170 => 170,
171 => 171,
172 => 172,
173 => 173,
174 => 174,
175 => 175,
176 => 176,
177 => 177,
178 => 178,
179 => 179,
180 => 180,
181 => 181,
182 => 182,
183 => 183,
184 => 184,
185 => 185,
186 => 186,
187 => 187,
188 => 188,
189 => 189,
190 => 190,
191 => 191,
192 => 192,
193 => 193,
194 => 194,
195 => 195,
196 => 196,
197 => 197,
198 => 198,
199 => 199,
200 => 200,
201 => 201,
202 => 202,
203 => 203,
204 => 204,
205 => 205,
206 => 206,
207 => 207,
208 => 208,
209 => 209,
210 => 210,
211 => 211,
212 => 212,
213 => 213,
214 => 214,
215 => 215,
216 => 216,
217 => 217,
218 => 218,
219 => 219,
220 => 220,
221 => 221,
222 => 222,
223 => 223,
224 => 224,
225 => 225,
226 => 226,
227 => 227,
228 => 228,
229 => 229,
230 => 230,
231 => 231,
232 => 232,
233 => 233,
234 => 234,
235 => 235,
236 => 236,
237 => 237,
238 => 238,
239 => 239,
240 => 240,
241 => 241,
242 => 242,
243 => 243,
244 => 244,
245 => 245,
246 => 246,
247 => 247,
248 => 248,
249 => 249,
250 => 250,
251 => 251,
252 => 252,
253 => 253,
254 => 254,
255 => 0,
256 => 1,
257 => 2,
258 => 3,
259 => 4,
260 => 5,
261 => 6,
262 => 7,
263 => 8,
264 => 9,
265 => 10,
266 => 11,
267 => 12,
268 => 13,
269 => 14,
270 => 15,
271 => 16,
272 => 17,
273 => 18,
274 => 19,
275 => 20,
276 => 21,
277 => 22,
278 => 23,
279 => 24,
280 => 25,
281 => 26,
282 => 27,
283 => 28,
284 => 29,
285 => 30,
286 => 31,
287 => 32,
288 => 33,
289 => 34,
290 => 35,
291 => 36,
292 => 37,
293 => 38,
294 => 39,
295 => 40,
296 => 41,
297 => 42,
298 => 43,
299 => 44,
300 => 45,
301 => 46,
302 => 47,
303 => 48,
304 => 49,
305 => 50,
306 => 51,
307 => 52,
308 => 53,
309 => 54,
310 => 55,
311 => 56,
312 => 57,
313 => 58,
314 => 59,
315 => 60,
316 => 61,
317 => 62,
318 => 63,
319 => 64,
320 => 65,
321 => 66,
322 => 67,
323 => 68,
324 => 69,
325 => 70,
326 => 71,
327 => 72,
328 => 73,
329 => 74,
330 => 75,
331 => 76,
332 => 77,
333 => 78,
334 => 79,
335 => 80,
336 => 81,
337 => 82,
338 => 83,
339 => 84,
340 => 85,
341 => 86,
342 => 87,
343 => 88,
344 => 89,
345 => 90,
346 => 91,
347 => 92,
348 => 93,
349 => 94,
350 => 95,
351 => 96,
352 => 97,
353 => 98,
354 => 99,
355 => 100,
356 => 101,
357 => 102,
358 => 103,
359 => 104,
360 => 105,
361 => 106,
362 => 107,
363 => 108,
364 => 109,
365 => 110,
366 => 111,
367 => 112,
368 => 113,
369 => 114,
370 => 115,
371 => 116,
372 => 117,
373 => 118,
374 => 119,
375 => 120,
376 => 121,
377 => 122,
378 => 123,
379 => 124,
380 => 125,
381 => 126,
382 => 127,
383 => 128,
384 => 129,
385 => 130,
386 => 131,
387 => 132,
388 => 133,
389 => 134,
390 => 135,
391 => 136,
392 => 137,
393 => 138,
394 => 139,
395 => 140,
396 => 141,
397 => 142,
398 => 143,
399 => 144,
400 => 145,
401 => 146,
402 => 147,
403 => 148,
404 => 149,
405 => 150,
406 => 151,
407 => 152,
408 => 153,
409 => 154,
410 => 155,
411 => 156,
412 => 157,
413 => 158,
414 => 159,
415 => 160,
416 => 161,
417 => 162,
418 => 163,
419 => 164,
420 => 165,
421 => 166,
422 => 167,
423 => 168,
424 => 169,
425 => 170,
426 => 171,
427 => 172,
428 => 173,
429 => 174,
430 => 175,
431 => 176,
432 => 177,
433 => 178,
434 => 179,
435 => 180,
436 => 181,
437 => 182,
438 => 183,
439 => 184,
440 => 185,
441 => 186,
442 => 187,
443 => 188,
444 => 189,
445 => 190,
446 => 191,
447 => 192,
448 => 193,
449 => 194,
450 => 195,
451 => 196,
452 => 197,
453 => 198,
454 => 199,
455 => 200,
456 => 201,
457 => 202,
458 => 203,
459 => 204,
460 => 205,
461 => 206,
462 => 207,
463 => 208,
464 => 209,
465 => 210,
466 => 211,
467 => 212,
468 => 213,
469 => 214,
470 => 215,
471 => 216,
472 => 217,
473 => 218,
474 => 219,
475 => 220,
476 => 221,
477 => 222,
478 => 223,
479 => 224,
480 => 225,
481 => 226,
482 => 227,
483 => 228,
484 => 229,
485 => 230,
486 => 231,
487 => 232,
488 => 233,
489 => 234,
490 => 235,
491 => 236,
492 => 237,
493 => 238,
494 => 239,
495 => 240,
496 => 241,
497 => 242,
498 => 243,
499 => 244,
500 => 245,
501 => 246,
502 => 247,
503 => 248,
504 => 249,
505 => 250,
506 => 251,
507 => 252,
508 => 253,
509 => 254,
510 => 0,
511 => 1,
512 => 2,
513 => 3,
514 => 4,
515 => 5,
516 => 6,
517 => 7,
518 => 8,
519 => 9,
520 => 10,
521 => 11,
522 => 12,
523 => 13,
524 => 14,
525 => 15,
526 => 16,
527 => 17,
528 => 18,
529 => 19,
530 => 20,
531 => 21,
532 => 22,
533 => 23,
534 => 24,
535 => 25,
536 => 26,
537 => 27,
538 => 28,
539 => 29,
540 => 30,
541 => 31,
542 => 32,
543 => 33,
544 => 34,
545 => 35,
546 => 36,
547 => 37,
548 => 38,
549 => 39,
550 => 40,
551 => 41,
552 => 42,
553 => 43,
554 => 44,
555 => 45,
556 => 46,
557 => 47,
558 => 48,
559 => 49,
560 => 50,
561 => 51,
562 => 52,
563 => 53,
564 => 54,
565 => 55,
566 => 56,
567 => 57,
568 => 58,
569 => 59,
570 => 60,
571 => 61,
572 => 62,
573 => 63,
574 => 64,
575 => 65,
576 => 66,
577 => 67,
578 => 68,
579 => 69,
580 => 70,
581 => 71,
582 => 72,
583 => 73,
584 => 74,
585 => 75,
586 => 76,
587 => 77,
588 => 78,
589 => 79,
590 => 80,
591 => 81,
592 => 82,
593 => 83,
594 => 84,
595 => 85,
596 => 86,
597 => 87,
598 => 88,
599 => 89,
600 => 90,
601 => 91,
602 => 92,
603 => 93,
604 => 94,
605 => 95,
606 => 96,
607 => 97,
608 => 98,
609 => 99,
610 => 100,
611 => 101,
612 => 102,
613 => 103,
614 => 104,
615 => 105,
616 => 106,
617 => 107,
618 => 108,
619 => 109,
620 => 110,
621 => 111,
622 => 112,
623 => 113,
624 => 114,
625 => 115,
626 => 116,
627 => 117,
628 => 118,
629 => 119,
630 => 120,
631 => 121,
632 => 122,
633 => 123,
634 => 124,
635 => 125,
636 => 126,
637 => 127,
638 => 128,
639 => 129,
640 => 130,
641 => 131,
642 => 132,
643 => 133,
644 => 134,
645 => 135,
646 => 136,
647 => 137,
648 => 138,
649 => 139,
650 => 140,
651 => 141,
652 => 142,
653 => 143,
654 => 144,
655 => 145,
656 => 146,
657 => 147,
658 => 148,
659 => 149,
660 => 150,
661 => 151,
662 => 152,
663 => 153,
664 => 154,
665 => 155,
666 => 156,
667 => 157,
668 => 158,
669 => 159,
670 => 160,
671 => 161,
672 => 162,
673 => 163,
674 => 164,
675 => 165,
676 => 166,
677 => 167,
678 => 168,
679 => 169,
680 => 170,
681 => 171,
682 => 172,
683 => 173,
684 => 174,
685 => 175,
686 => 176,
687 => 177,
688 => 178,
689 => 179,
690 => 180,
691 => 181,
692 => 182,
693 => 183,
694 => 184,
695 => 185,
696 => 186,
697 => 187,
698 => 188,
699 => 189,
700 => 190,
701 => 191,
702 => 192,
703 => 193,
704 => 194,
705 => 195,
706 => 196,
707 => 197,
708 => 198,
709 => 199,
710 => 200,
711 => 201,
712 => 202,
713 => 203,
714 => 204,
715 => 205,
716 => 206,
717 => 207,
718 => 208,
719 => 209,
720 => 210,
721 => 211,
722 => 212,
723 => 213,
724 => 214,
725 => 215,
726 => 216,
727 => 217,
728 => 218,
729 => 219,
730 => 220,
731 => 221,
732 => 222,
733 => 223,
734 => 224,
735 => 225,
736 => 226,
737 => 227,
738 => 228,
739 => 229,
740 => 230,
741 => 231,
742 => 232,
743 => 233,
744 => 234,
745 => 235,
746 => 236,
747 => 237,
748 => 238,
749 => 239,
750 => 240,
751 => 241,
752 => 242,
753 => 243,
754 => 244,
755 => 245,
756 => 246,
757 => 247,
758 => 248,
759 => 249,
760 => 250,
761 => 251,
762 => 252,
763 => 253,
764 => 254,
765 => 0
);

signal test, outputtemp, epattern1, epattern2, epattern : std_logic_vector(254 downto 0);
signal S1 : std_logic_vector(7 downto 0);
signal S3 : std_logic_vector(7 downto 0);
signal s1pow3, s3pow1, s1pow3s3 : integer;
signal rat : std_logic_vector(7 downto 0);
signal y1, y2, e1pos, e2pos : integer range 0 to 255;

component Syndrome1Calc is
	port( 
		R  : in std_logic_vector(254 downto 0); 
		output : out std_logic_vector(7 downto 0)
	);
end component;

component Syndrome3Calc is
	port( 
		R  : in std_logic_vector(254 downto 0); 
		output : out std_logic_vector(7 downto 0)
	);
end component;

begin


--S1 as exponent of primitive element to the third power
--polyval(S1, 2)

process(clock,input)
begin
--test <= "111000110010101000000110100001100100000010000111110110111110000110110010101011100010001110000010010001100000000101101110000101000111010001110100011101010100001011100101101111001000101010001111101010100011011100011000101100001010111110110100100101110011011";
test <= input;
end process;

process (S1, clock)
begin
	if (to_integer(unsigned(S1)) > 0) then
		s1pow3 <= ROM_MOD(ROM_alphaInv(to_integer(unsigned(S1)))*3); --log(s1^3)
  end if;
end process;

--% S3 as exponent of primitive element
process (S3)
begin
	if (to_integer(unsigned(S3)) > 0) then
		s3pow1 <= ROM_alphaInv(to_integer(unsigned(S3))); --log(s3)
  end if;
end process;


--% Subtracting the exponents 
--A = sigma2 / sigma1^2
s1pow3s3 <= ROM_MOD((s3pow1 - s1pow3));


process (s1pow3s3, S3) --rat = bitxor(alpha(s1pow3s3+1,:), alpha(0+1,:));
begin
	if (s1pow3s3 >= 0) then
	
		if (S3 = "00000000") then
			rat <= ROM_alpha(1);
		else
			rat <= ROM_alpha((s1pow3s3+1)) xor ROM_alpha(1);
		end if;
	
	end if;
end process;


process(rat)
begin
if (to_integer(unsigned(rat)) > 0) then
y1 <= ROM_yFirstMatch(ROM_alphaInv(to_integer(unsigned(rat))));
y2 <= ROM_ySecondMatch(ROM_alphaInv(to_integer(unsigned(rat))));
end if;
end process;


process(y1,y2,clock) --x = 255 - mod(y+alphainv(BinToDec(S1),:), 2^m - 1);
begin

if (to_integer(unsigned(S1)) > 0) then --- MINUS 1 because of the VHLD indexing
e1pos <= (255 - (ROM_MOD(y1 + ROM_alphaInv(to_integer(unsigned(S1))) ))) -1;
e2pos <= (255 - (ROM_MOD(y2 + ROM_alphaInv(to_integer(unsigned(S1))) ))) -1;
end if;

end process;


process(e1pos,e2pos) --x = 255 - mod(y+alphainv(BinToDec(S1),:), 2^m - 1);
begin

if (y1 > 0 or y2 > 0) then
epattern1 <= ROM_E(e1pos+1);
epattern2 <= ROM_E(e2pos+1);
--epattern1 <= (e1pos      => '1',
--			  others => '0');
--epattern2 <= (e2pos      => '1',
--			  others => '0');
else
epattern1 <= ROM_E(0);
epattern2 <= ROM_E(0);

end if;

end process;


process(epattern1,epattern2) --x = 255 - mod(y+alphainv(BinToDec(S1),:), 2^m - 1);
begin

epattern <= epattern1 xor epattern2;

outputtemp <= test;

end process;

process(epattern) --x = 255 - mod(y+alphainv(BinToDec(S1),:), 2^m - 1);
begin

output <= epattern xor outputtemp;

end process;

DUT1 : Syndrome1Calc
	port map(
		R  => test,
		output => S1
	);

DUT2 : Syndrome3Calc
	port map(
		R  => test,
		output => S3
	);

end architecture;


