LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

entity Syndrome1Calc is
	port( 
		R  : in std_logic_vector(254 downto 0); 
		output : out std_logic_vector(7 downto 0)
	);
end entity;

architecture Syndrome1Calc_arch of Syndrome1Calc is

signal S1 : std_logic_vector(7 downto 0);

begin

S1(0) <= R(0) xor R(2) xor R(3) xor R(7) xor R(8) xor R(9) xor R(10) xor R(12) xor R(17) xor R(18) xor R(19) xor R(20) xor R(21) xor R(22) xor R(23) xor R(24) xor R(27) xor R(32) xor R(34) xor R(37) xor R(38) xor R(39) xor R(40) xor R(41) xor R(43) xor R(45) xor R(47) xor R(49) xor R(50) xor R(51) xor R(57) xor R(58) xor R(62) xor R(64) xor R(66) xor R(67) xor R(70) xor R(71) xor R(74) xor R(76) xor R(77) xor R(78) xor R(79) xor R(80) xor R(81) xor R(83) xor R(84) xor R(85) xor R(86) xor R(89) xor R(90) xor R(92) xor R(93) xor R(94) xor R(96) xor R(97) xor R(98) xor R(101) xor R(103) xor R(105) xor R(108) xor R(110) xor R(114) xor R(117) xor R(119) xor R(120) xor R(122) xor R(126) xor R(127) xor R(130) xor R(131) xor R(132) xor R(135) xor R(136) xor R(137) xor R(138) xor R(142) xor R(143) xor R(145) xor R(146) xor R(151) xor R(155) xor R(157) xor R(158) xor R(159) xor R(161) xor R(163) xor R(164) xor R(165) xor R(166) xor R(168) xor R(169) xor R(171) xor R(172) xor R(173) xor R(174) xor R(175) xor R(180) xor R(181) xor R(183) xor R(186) xor R(187) xor R(189) xor R(191) xor R(192) xor R(194) xor R(195) xor R(197) xor R(199) xor R(205) xor R(208) xor R(209) xor R(210) xor R(212) xor R(213) xor R(216) xor R(219) xor R(222) xor R(223) xor R(230) xor R(231) xor R(232) xor R(234) xor R(237) xor R(241) xor R(242) xor R(243) xor R(247) ;
S1(1) <= R(1) xor R(3) xor R(4) xor R(8) xor R(9) xor R(10) xor R(11) xor R(13) xor R(18) xor R(19) xor R(20) xor R(21) xor R(22) xor R(23) xor R(24) xor R(25) xor R(28) xor R(33) xor R(35) xor R(38) xor R(39) xor R(40) xor R(41) xor R(42) xor R(44) xor R(46) xor R(48) xor R(50) xor R(51) xor R(52) xor R(58) xor R(59) xor R(63) xor R(65) xor R(67) xor R(68) xor R(71) xor R(72) xor R(75) xor R(77) xor R(78) xor R(79) xor R(80) xor R(81) xor R(82) xor R(84) xor R(85) xor R(86) xor R(87) xor R(90) xor R(91) xor R(93) xor R(94) xor R(95) xor R(97) xor R(98) xor R(99) xor R(102) xor R(104) xor R(106) xor R(109) xor R(111) xor R(115) xor R(118) xor R(120) xor R(121) xor R(123) xor R(127) xor R(128) xor R(131) xor R(132) xor R(133) xor R(136) xor R(137) xor R(138) xor R(139) xor R(143) xor R(144) xor R(146) xor R(147) xor R(152) xor R(156) xor R(158) xor R(159) xor R(160) xor R(162) xor R(164) xor R(165) xor R(166) xor R(167) xor R(169) xor R(170) xor R(172) xor R(173) xor R(174) xor R(175) xor R(176) xor R(181) xor R(182) xor R(184) xor R(187) xor R(188) xor R(190) xor R(192) xor R(193) xor R(195) xor R(196) xor R(198) xor R(200) xor R(206) xor R(209) xor R(210) xor R(211) xor R(213) xor R(214) xor R(217) xor R(220) xor R(223) xor R(224) xor R(231) xor R(232) xor R(233) xor R(235) xor R(238) xor R(242) xor R(243) xor R(244) xor R(248) ;
S1(2) <= R(2) xor R(4) xor R(5) xor R(9) xor R(10) xor R(11) xor R(12) xor R(14) xor R(19) xor R(20) xor R(21) xor R(22) xor R(23) xor R(24) xor R(25) xor R(26) xor R(29) xor R(34) xor R(36) xor R(39) xor R(40) xor R(41) xor R(42) xor R(43) xor R(45) xor R(47) xor R(49) xor R(51) xor R(52) xor R(53) xor R(59) xor R(60) xor R(64) xor R(66) xor R(68) xor R(69) xor R(72) xor R(73) xor R(76) xor R(78) xor R(79) xor R(80) xor R(81) xor R(82) xor R(83) xor R(85) xor R(86) xor R(87) xor R(88) xor R(91) xor R(92) xor R(94) xor R(95) xor R(96) xor R(98) xor R(99) xor R(100) xor R(103) xor R(105) xor R(107) xor R(110) xor R(112) xor R(116) xor R(119) xor R(121) xor R(122) xor R(124) xor R(128) xor R(129) xor R(132) xor R(133) xor R(134) xor R(137) xor R(138) xor R(139) xor R(140) xor R(144) xor R(145) xor R(147) xor R(148) xor R(153) xor R(157) xor R(159) xor R(160) xor R(161) xor R(163) xor R(165) xor R(166) xor R(167) xor R(168) xor R(170) xor R(171) xor R(173) xor R(174) xor R(175) xor R(176) xor R(177) xor R(182) xor R(183) xor R(185) xor R(188) xor R(189) xor R(191) xor R(193) xor R(194) xor R(196) xor R(197) xor R(199) xor R(201) xor R(207) xor R(210) xor R(211) xor R(212) xor R(214) xor R(215) xor R(218) xor R(221) xor R(224) xor R(225) xor R(232) xor R(233) xor R(234) xor R(236) xor R(239) xor R(243) xor R(244) xor R(245) xor R(249) ;
S1(3) <= R(3) xor R(5) xor R(6) xor R(10) xor R(11) xor R(12) xor R(13) xor R(15) xor R(20) xor R(21) xor R(22) xor R(23) xor R(24) xor R(25) xor R(26) xor R(27) xor R(30) xor R(35) xor R(37) xor R(40) xor R(41) xor R(42) xor R(43) xor R(44) xor R(46) xor R(48) xor R(50) xor R(52) xor R(53) xor R(54) xor R(60) xor R(61) xor R(65) xor R(67) xor R(69) xor R(70) xor R(73) xor R(74) xor R(77) xor R(79) xor R(80) xor R(81) xor R(82) xor R(83) xor R(84) xor R(86) xor R(87) xor R(88) xor R(89) xor R(92) xor R(93) xor R(95) xor R(96) xor R(97) xor R(99) xor R(100) xor R(101) xor R(104) xor R(106) xor R(108) xor R(111) xor R(113) xor R(117) xor R(120) xor R(122) xor R(123) xor R(125) xor R(129) xor R(130) xor R(133) xor R(134) xor R(135) xor R(138) xor R(139) xor R(140) xor R(141) xor R(145) xor R(146) xor R(148) xor R(149) xor R(154) xor R(158) xor R(160) xor R(161) xor R(162) xor R(164) xor R(166) xor R(167) xor R(168) xor R(169) xor R(171) xor R(172) xor R(174) xor R(175) xor R(176) xor R(177) xor R(178) xor R(183) xor R(184) xor R(186) xor R(189) xor R(190) xor R(192) xor R(194) xor R(195) xor R(197) xor R(198) xor R(200) xor R(202) xor R(208) xor R(211) xor R(212) xor R(213) xor R(215) xor R(216) xor R(219) xor R(222) xor R(225) xor R(226) xor R(233) xor R(234) xor R(235) xor R(237) xor R(240) xor R(244) xor R(245) xor R(246) xor R(250) ;
S1(4) <= R(0) xor R(2) xor R(3) xor R(4) xor R(6) xor R(8) xor R(9) xor R(10) xor R(11) xor R(13) xor R(14) xor R(16) xor R(17) xor R(18) xor R(19) xor R(20) xor R(25) xor R(26) xor R(28) xor R(31) xor R(32) xor R(34) xor R(36) xor R(37) xor R(39) xor R(40) xor R(42) xor R(44) xor R(50) xor R(53) xor R(54) xor R(55) xor R(57) xor R(58) xor R(61) xor R(64) xor R(67) xor R(68) xor R(75) xor R(76) xor R(77) xor R(79) xor R(82) xor R(86) xor R(87) xor R(88) xor R(92) xor R(100) xor R(102) xor R(103) xor R(107) xor R(108) xor R(109) xor R(110) xor R(112) xor R(117) xor R(118) xor R(119) xor R(120) xor R(121) xor R(122) xor R(123) xor R(124) xor R(127) xor R(132) xor R(134) xor R(137) xor R(138) xor R(139) xor R(140) xor R(141) xor R(143) xor R(145) xor R(147) xor R(149) xor R(150) xor R(151) xor R(157) xor R(158) xor R(162) xor R(164) xor R(166) xor R(167) xor R(170) xor R(171) xor R(174) xor R(176) xor R(177) xor R(178) xor R(179) xor R(180) xor R(181) xor R(183) xor R(184) xor R(185) xor R(186) xor R(189) xor R(190) xor R(192) xor R(193) xor R(194) xor R(196) xor R(197) xor R(198) xor R(201) xor R(203) xor R(205) xor R(208) xor R(210) xor R(214) xor R(217) xor R(219) xor R(220) xor R(222) xor R(226) xor R(227) xor R(230) xor R(231) xor R(232) xor R(235) xor R(236) xor R(237) xor R(238) xor R(242) xor R(243) xor R(245) xor R(246) xor R(251) ;
S1(5) <= R(0) xor R(1) xor R(2) xor R(4) xor R(5) xor R(8) xor R(11) xor R(14) xor R(15) xor R(22) xor R(23) xor R(24) xor R(26) xor R(29) xor R(33) xor R(34) xor R(35) xor R(39) xor R(47) xor R(49) xor R(50) xor R(54) xor R(55) xor R(56) xor R(57) xor R(59) xor R(64) xor R(65) xor R(66) xor R(67) xor R(68) xor R(69) xor R(70) xor R(71) xor R(74) xor R(79) xor R(81) xor R(84) xor R(85) xor R(86) xor R(87) xor R(88) xor R(90) xor R(92) xor R(94) xor R(96) xor R(97) xor R(98) xor R(104) xor R(105) xor R(109) xor R(111) xor R(113) xor R(114) xor R(117) xor R(118) xor R(121) xor R(123) xor R(124) xor R(125) xor R(126) xor R(127) xor R(128) xor R(130) xor R(131) xor R(132) xor R(133) xor R(136) xor R(137) xor R(139) xor R(140) xor R(141) xor R(143) xor R(144) xor R(145) xor R(148) xor R(150) xor R(152) xor R(155) xor R(157) xor R(161) xor R(164) xor R(166) xor R(167) xor R(169) xor R(173) xor R(174) xor R(177) xor R(178) xor R(179) xor R(182) xor R(183) xor R(184) xor R(185) xor R(189) xor R(190) xor R(192) xor R(193) xor R(198) xor R(202) xor R(204) xor R(205) xor R(206) xor R(208) xor R(210) xor R(211) xor R(212) xor R(213) xor R(215) xor R(216) xor R(218) xor R(219) xor R(220) xor R(221) xor R(222) xor R(227) xor R(228) xor R(230) xor R(233) xor R(234) xor R(236) xor R(238) xor R(239) xor R(241) xor R(242) xor R(244) xor R(246) xor R(252) ;
S1(6) <= R(0) xor R(1) xor R(5) xor R(6) xor R(7) xor R(8) xor R(10) xor R(15) xor R(16) xor R(17) xor R(18) xor R(19) xor R(20) xor R(21) xor R(22) xor R(25) xor R(30) xor R(32) xor R(35) xor R(36) xor R(37) xor R(38) xor R(39) xor R(41) xor R(43) xor R(45) xor R(47) xor R(48) xor R(49) xor R(55) xor R(56) xor R(60) xor R(62) xor R(64) xor R(65) xor R(68) xor R(69) xor R(72) xor R(74) xor R(75) xor R(76) xor R(77) xor R(78) xor R(79) xor R(81) xor R(82) xor R(83) xor R(84) xor R(87) xor R(88) xor R(90) xor R(91) xor R(92) xor R(94) xor R(95) xor R(96) xor R(99) xor R(101) xor R(103) xor R(106) xor R(108) xor R(112) xor R(115) xor R(117) xor R(118) xor R(120) xor R(124) xor R(125) xor R(128) xor R(129) xor R(130) xor R(133) xor R(134) xor R(135) xor R(136) xor R(140) xor R(141) xor R(143) xor R(144) xor R(149) xor R(153) xor R(155) xor R(156) xor R(157) xor R(159) xor R(161) xor R(162) xor R(163) xor R(164) xor R(166) xor R(167) xor R(169) xor R(170) xor R(171) xor R(172) xor R(173) xor R(178) xor R(179) xor R(181) xor R(184) xor R(185) xor R(187) xor R(189) xor R(190) xor R(192) xor R(193) xor R(195) xor R(197) xor R(203) xor R(206) xor R(207) xor R(208) xor R(210) xor R(211) xor R(214) xor R(217) xor R(220) xor R(221) xor R(228) xor R(229) xor R(230) xor R(232) xor R(235) xor R(239) xor R(240) xor R(241) xor R(245) xor R(253) ;
S1(7) <= R(1) xor R(2) xor R(6) xor R(7) xor R(8) xor R(9) xor R(11) xor R(16) xor R(17) xor R(18) xor R(19) xor R(20) xor R(21) xor R(22) xor R(23) xor R(26) xor R(31) xor R(33) xor R(36) xor R(37) xor R(38) xor R(39) xor R(40) xor R(42) xor R(44) xor R(46) xor R(48) xor R(49) xor R(50) xor R(56) xor R(57) xor R(61) xor R(63) xor R(65) xor R(66) xor R(69) xor R(70) xor R(73) xor R(75) xor R(76) xor R(77) xor R(78) xor R(79) xor R(80) xor R(82) xor R(83) xor R(84) xor R(85) xor R(88) xor R(89) xor R(91) xor R(92) xor R(93) xor R(95) xor R(96) xor R(97) xor R(100) xor R(102) xor R(104) xor R(107) xor R(109) xor R(113) xor R(116) xor R(118) xor R(119) xor R(121) xor R(125) xor R(126) xor R(129) xor R(130) xor R(131) xor R(134) xor R(135) xor R(136) xor R(137) xor R(141) xor R(142) xor R(144) xor R(145) xor R(150) xor R(154) xor R(156) xor R(157) xor R(158) xor R(160) xor R(162) xor R(163) xor R(164) xor R(165) xor R(167) xor R(168) xor R(170) xor R(171) xor R(172) xor R(173) xor R(174) xor R(179) xor R(180) xor R(182) xor R(185) xor R(186) xor R(188) xor R(190) xor R(191) xor R(193) xor R(194) xor R(196) xor R(198) xor R(204) xor R(207) xor R(208) xor R(209) xor R(211) xor R(212) xor R(215) xor R(218) xor R(221) xor R(222) xor R(229) xor R(230) xor R(231) xor R(233) xor R(236) xor R(240) xor R(241) xor R(242) xor R(246) xor R(254) ;

output <= S1;
	
end architecture;
