
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

entity test is
end entity;

architecture test_arch of test is

signal testvektor : std_logic_vector(3 downto 0);
signal umm : std_logic_vector(3 downto 0);

type ROM_type is array (0 to 254) of std_logic_vector(7 downto 0);
constant ROM_alpha : ROM_type := ( 0 => "00000001",
1 => "00000010",
2 => "00000100",
3 => "00001000",
4 => "00010000",
5 => "00100000",
6 => "01000000",
7 => "10000000",
8 => "00011101",
9 => "00111010",
10 => "01110100",
11 => "11101000",
12 => "11001101",
13 => "10000111",
14 => "00010011",
15 => "00100110",
16 => "01001100",
17 => "10011000",
18 => "00101101",
19 => "01011010",
20 => "10110100",
21 => "01110101",
22 => "11101010",
23 => "11001001",
24 => "10001111",
25 => "00000011",
26 => "00000110",
27 => "00001100",
28 => "00011000",
29 => "00110000",
30 => "01100000",
31 => "11000000",
32 => "10011101",
33 => "00100111",
34 => "01001110",
35 => "10011100",
36 => "00100101",
37 => "01001010",
38 => "10010100",
39 => "00110101",
40 => "01101010",
41 => "11010100",
42 => "10110101",
43 => "01110111",
44 => "11101110",
45 => "11000001",
46 => "10011111",
47 => "00100011",
48 => "01000110",
49 => "10001100",
50 => "00000101",
51 => "00001010",
52 => "00010100",
53 => "00101000",
54 => "01010000",
55 => "10100000",
56 => "01011101",
57 => "10111010",
58 => "01101001",
59 => "11010010",
60 => "10111001",
61 => "01101111",
62 => "11011110",
63 => "10100001",
64 => "01011111",
65 => "10111110",
66 => "01100001",
67 => "11000010",
68 => "10011001",
69 => "00101111",
70 => "01011110",
71 => "10111100",
72 => "01100101",
73 => "11001010",
74 => "10001001",
75 => "00001111",
76 => "00011110",
77 => "00111100",
78 => "01111000",
79 => "11110000",
80 => "11111101",
81 => "11100111",
82 => "11010011",
83 => "10111011",
84 => "01101011",
85 => "11010110",
86 => "10110001",
87 => "01111111",
88 => "11111110",
89 => "11100001",
90 => "11011111",
91 => "10100011",
92 => "01011011",
93 => "10110110",
94 => "01110001",
95 => "11100010",
96 => "11011001",
97 => "10101111",
98 => "01000011",
99 => "10000110",
100 => "00010001",
101 => "00100010",
102 => "01000100",
103 => "10001000",
104 => "00001101",
105 => "00011010",
106 => "00110100",
107 => "01101000",
108 => "11010000",
109 => "10111101",
110 => "01100111",
111 => "11001110",
112 => "10000001",
113 => "00011111",
114 => "00111110",
115 => "01111100",
116 => "11111000",
117 => "11101101",
118 => "11000111",
119 => "10010011",
120 => "00111011",
121 => "01110110",
122 => "11101100",
123 => "11000101",
124 => "10010111",
125 => "00110011",
126 => "01100110",
127 => "11001100",
128 => "10000101",
129 => "00010111",
130 => "00101110",
131 => "01011100",
132 => "10111000",
133 => "01101101",
134 => "11011010",
135 => "10101001",
136 => "01001111",
137 => "10011110",
138 => "00100001",
139 => "01000010",
140 => "10000100",
141 => "00010101",
142 => "00101010",
143 => "01010100",
144 => "10101000",
145 => "01001101",
146 => "10011010",
147 => "00101001",
148 => "01010010",
149 => "10100100",
150 => "01010101",
151 => "10101010",
152 => "01001001",
153 => "10010010",
154 => "00111001",
155 => "01110010",
156 => "11100100",
157 => "11010101",
158 => "10110111",
159 => "01110011",
160 => "11100110",
161 => "11010001",
162 => "10111111",
163 => "01100011",
164 => "11000110",
165 => "10010001",
166 => "00111111",
167 => "01111110",
168 => "11111100",
169 => "11100101",
170 => "11010111",
171 => "10110011",
172 => "01111011",
173 => "11110110",
174 => "11110001",
175 => "11111111",
176 => "11100011",
177 => "11011011",
178 => "10101011",
179 => "01001011",
180 => "10010110",
181 => "00110001",
182 => "01100010",
183 => "11000100",
184 => "10010101",
185 => "00110111",
186 => "01101110",
187 => "11011100",
188 => "10100101",
189 => "01010111",
190 => "10101110",
191 => "01000001",
192 => "10000010",
193 => "00011001",
194 => "00110010",
195 => "01100100",
196 => "11001000",
197 => "10001101",
198 => "00000111",
199 => "00001110",
200 => "00011100",
201 => "00111000",
202 => "01110000",
203 => "11100000",
204 => "11011101",
205 => "10100111",
206 => "01010011",
207 => "10100110",
208 => "01010001",
209 => "10100010",
210 => "01011001",
211 => "10110010",
212 => "01111001",
213 => "11110010",
214 => "11111001",
215 => "11101111",
216 => "11000011",
217 => "10011011",
218 => "00101011",
219 => "01010110",
220 => "10101100",
221 => "01000101",
222 => "10001010",
223 => "00001001",
224 => "00010010",
225 => "00100100",
226 => "01001000",
227 => "10010000",
228 => "00111101",
229 => "01111010",
230 => "11110100",
231 => "11110101",
232 => "11110111",
233 => "11110011",
234 => "11111011",
235 => "11101011",
236 => "11001011",
237 => "10001011",
238 => "00001011",
239 => "00010110",
240 => "00101100",
241 => "01011000",
242 => "10110000",
243 => "01111101",
244 => "11111010",
245 => "11101001",
246 => "11001111",
247 => "10000011",
248 => "00011011",
249 => "00110110",
250 => "01101100",
251 => "11011000",
252 => "10101101",
253 => "01000111",
254 => "10001110"
);

begin
	
umm <= "0011";
	
testvektor(0) <= '0' xor umm(0);
testvektor(1) <= '1' xor umm(1);
testvektor(2) <= '0' xor umm(2);
testvektor(3) <= '1' xor umm(3);



end architecture;
