LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
USE IEEE.std_logic_textio.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

LIBRARY STD;
USE STD.textio.all;

entity Decoder_TB is
end entity;

architecture Decoder_TB_arch of Decoder_TB is

component Decoder is
		port(  
		clock  : in std_logic;
		input  : std_logic_vector(254 downto 0);
		output : out std_logic_vector(254 downto 0)
		);
end component;

--TB clock
signal Clock, ok : std_logic;
constant clk_period: time:=10 ns;
signal result : std_logic_vector(254 downto 0);
signal test, check  : std_logic_vector(254 downto 0);
signal counter : integer range 1 to 100;

--FOR SINGLE TESTING
type ROM_typeSingle is array (0 to 0) of std_logic_vector(254 downto 0);
constant ROM_SINGLEin : ROM_typeSingle := ( 
0 =>  "000001001100101001011110101101011011010010100100111001110001101000001001101010000010011100000100010010011101111101001110100010110011111110100110111010001101110010001100010010011100011111000111100110010110011010111010100011110010100101011101101110000010100"
);
constant ROM_SINGLEout : ROM_typeSingle := ( 
0 => "000001001100101001011010101101011011010010100100111001111001101000001001101010000010011100000100010010011101111101001110100010110011111110100110111010001101110010001100010010011100011111000111100110010110011010111010100011110010100101011101101110000010100"
);


--000001001100101001011110101101011011010010100100111001110001101000001001101010000010011100000100010010011101111101001110100010110011111110100110111010001101110010001100010010011100011111000111100110010110011010111010100011110010100101011101101110000010100
--000001001100101001011810101101011011010010100100111001118001101000001001101010000010011100000100010010011101111101001110100010110011111110100110111010001101110010001100010010011100011111000111100110010110011010111010100011110010100101011101101110000010100
--


type ROM_type is array (1 to 100) of std_logic_vector(254 downto 0);
constant ROM_C : ROM_type := ( 1 => "101101101010001000101000000101101000010001011010110010000100001000010101111011110000000101010001000011101010101011101000100111111000100101000100000110110000000110110010110110110100000000010011001001000010001010011000010011110100001110001011001100101111101",
2 => "010011111110011100101000101011111010001101110000110001000001111100010011111000000100011111101110000010001010110111011000110010111001111110110000111011101100100001011101111110110011001000011010111101100100110110001011100010100101100000110101011101011011010",
3 => "010000000110100101111010010000000011001100010110101000110110011011011111100001110111111100001110001010010001000001000000011000011001101011001000000001101111111000010010101001100110011100011110010001110110011101101001111000110000101110001111111000110111110",
4 => "011010011111001010111000110100001111100011110000001100001111101010001101001110111110100111111000111001111100110000010011000110111110010111111001000000100100011111111000010010001010101001100001110101111010111111101000101011101111010111101000010110110111101",
5 => "101101000010000110010110000000110001001000110101010110101000100110111100111011010110101100100111011000100100111111100010111100110111100110001011001101000001100011110000100101011001010101000010000000110110001101101000000011111000010101111010110111110110101",
6 => "001000100001110110011110101100110001110101110010000101010011100110111010110001000111001011100001101010011101101000111000001001111111000010100000000111000111111000111011101100101000111000111110100111111101101010100010100001000000000110010000110110011011101",
7 => "101111010010101000111010110111100111001111001111010101011101100011001101100101000111011101000011111000110100010001000011010010110101010100010111000110000111010010101001101010110001010000000010000101010010100101000011011010110100000110100010000101011000011",
8 => "010000011001000100000101011101110110001011101111110000010011110111110100011110001010010000111000111110101100000101011000100000101100111001000111110100110010101100001010101101101101000001000101110000010000101100101000001011011001011001101101011110110000010",
9 => "101000011101000101011111000001001011011010010110100001011101101001010101011011110010101001001101101001111001001110100000001100101100111100011111101111111100011000101110011100011100000011011001000111010100010111111100000001100011001110010000010001100111001",
10 => "100110111110101101001111011011000110000000101011011001000000100100111111001000101010011101100011010111101000000111111101101100011010101011111000001001010110010101010101111011111001101000111010100111111100101100101011101011101111101111111110111001001111101",
11 => "110010101001001000100100110001110001011110001111100011000010100100010100000000110110011001101001100011111010000111011100011011101111111000111001001100011110010001100111100000001100111001000001000000011110110011100010100000001101111010101010101010001000000",
12 => "110010000001110001001010101011100001110111111010111010101011111110010100010101111001011011010011011000111010100001110011100011001001000000110110000110011101110100000001001000101100011001011100010000111001101111111111110101011100001111011110111010011100101",
13 => "011011000110100011101011100000000111000000100010010001110010100000010110000001101101101101011111010110101010100110110110011011010101110110011111110000101110001101110001011011011101110100010110010010000110100011000011100110011001111101001100111001101011111",
14 => "010101101001110010101000011101110011110011110100010100011001010110101101111011001100010100100110010101111000110000001001100100000101110010101001111001011111100011010111111111100100111001001101100110110000000000001011011110000001100101000000010101111111100",
15 => "110100011111100010000111101111001001000001111100111101110110100111001011001001011000000001000111011100111011100100000000111100101001000011000001101100111101011100010000101010111001001100111001110000101110010100010000010111101001111000101100101100000010001",
16 => "110011100000001010110000100000000011100010011111001111101010100101111111101001110101000000011101111101000000100011010100111110111110101010000001000111111010001100111000010100010100010001101000101000111011110001111110001000101011101111111001101111010010111",
17 => "110000010111011100000111100000001001111100000111111000011001110101101111111100011100100010100100010101101110010101001010110011011000111101101111000110100111101010110111100000001101011111110000110101001111000001000011110011111110101111001010000001010001000",
18 => "010110100000110011010111101000010001100101001111100010110000010110100001010110000110001111011111001000110000111101110011101111101110111001001100000011001101001111101000000000111111111110101000011011000111011000011000101110111000101001111111100111010000011",
19 => "001010000100001110111011110101101101000000100001100010110010101000000011011000001111100110100101010100111100000100010111101100111000101010011111111111111110010000011001100011001010000011100101000100110111101100010011111001000010111000110100110000000011111",
20 => "000010110101101000111110100001000011001000111010000111111010100011011110110100001010110001001001010111110111100100101001001100111010001010110011001010011111000010101010111101000001110010100000111010100111010100101101011000101011001010000001000111111101111",
21 => "010000101000100101110100111011001001011100110000011010000100110011001001001111011100111011010110000010010010100100010101000111100010001001011111010010100100011011101110110100101110000001110100111110001001011001011101110111010010011000110011100000001010001",
22 => "011100001000111111011101010111111100010110110010111001011011101101111011001101000101001011101111001110001010101011010111111110001010010100000110001011011011111110010010100111011010011100011001011001101001110010010101011001100111101101000110100000011100011",
23 => "111111101100110101001101001010010000010011100001100100110100101100000010011111100100110111101001111100000101100011010101111101110110011110000010010101001000100110011111011101010000001001111110101100001010000100001110100111100001101000010110000110010100100",
24 => "100011110110111110011001101010011011110000010111111001011011000110010111101010100001111100111100111000001100100110101001001010101101100000101110000111010101111001001010101010111000101010001111110011101001100010111100110010011110010101100101110110001110100",
25 => "011101001010100111110001100001111110100010010011101001010101010100010011010001111001001000110100111011110101010101011100010001000011101000110111010001000101111001000000001011100101000110000101010111001111101001110101101011001101000110000010011100110010110",
26 => "100010100101001000001001010100011100001111011010111001011000110101111101000010001111010101110100011100111110001111111001001000101111111110010100100001111010010001001001110101110110101100111011101100111110000100101011110111011100111101000010000111111101010",
27 => "100001011110000010100010111110100110011101111100001100110101100101101001000101101101001101010101110111001011011101001110110010101101100100010011100111010000010000000101100110000101111011010101111000010110001111000000100000000010000101111111010011001010011",
28 => "010011011010001100010110011110101011100000101011100100111110010000111011110111001011001010101110111011011100101111010011101011011110010111100000110100000000110100100001111101011101100001111110101011011100000001000000101001001101110010100011101001101010111",
29 => "000110100101110011111110011110110010111001111111100110101100010100000010010101100110101110011011110110011011100111101101111000000100001111000011101111000110110101110000000010000101000011100101000010010100100001011101100000010000101001101011011100111011110",
30 => "011010100110101010100010010101101000000110101111100001000111111001001011011011011001100101110100101001011110101000001110101101001111100111111000010101001001010110011000000000001011001100101010011010010001101000100000100110101111110101100100101010100101001",
31 => "101111111110100100011010000011000101100001001101100110100101000011001000101100111010100000001111001010100101010010001100000000001000011001100110111010100001111001011010010010111110000110111001010011001000001000011110100010100010000010101111000110110001100",
32 => "010101101001011101010100001010111010100001100000000001001101100100111111100001011011010111001000111011111001101010001111001000000110101000100000010010111101101011000011001101001001001001001101000111010001110101001000110110110110111010000011110101111100001",
33 => "110100011111000010100011110111001000000010000010110110011100000110111000001000101000001010011001001100111010110010100101010100001101000101011000100101010011010110111110000101001100001100011010000100110100100010000101000101100100101011110100010101110000001",
34 => "010011111000001010001001000110111011111110110010000001110011111110100000010010101001011000110001111100010001000110001011100001111110100111010110010100101101001100111000101111111001001110101001110110001110111110100111110011100011111000101001010110100101001",
35 => "100111110111001110000000011111101010000111110100001000011111110100100000100111000001100110110000011011010001100111011011101000101011101010100100111001010111000110100001000011111011101000100101000000010100000111101001000001001000110111001110110011001101111",
36 => "000000001000101011001001111101001011101000110000000110110101101100110010001011101001111000000110111110101010110100100011111010010101000101010010001101110101111111110111110100001000000010010001010000111110000100110110000101111111000001100000101001001010100",
37 => "001100100101111110111010001010011010110011000010011001000100011100001111001001110110100101011100000000110111011101101101101110100011100010001101111101011011010001100100000111010010110010101010011101010011011000010111100010010101100001100110101011010001010",
38 => "111010011110011010101001101010011001100000111001100100111010100010001011110000001010010100111111111000111010001100011110000111101011100100010000000101000110011100010001010100111111001000101111011111101011001100110011001101100000011101011011001111001001111",
39 => "100000011110010101010110100001010110011011100011010011010110100001010001011101110100010010010111100111110101010101011010010111001101111001000110101100100110000001000101010011010010010111110101010011011001111100001011101001100100110111001010011000000000000",
40 => "111100100111001001010000011101011010000111110010000101001011100110110101111100111000100101101001010110001111110001110000000100001001010110100101000100110010101110100010000000000000101011101101111110101001001111000010101011110111011001010001111000100011001",
41 => "001101110101010100001011000100001101100101111101011000000010111110001101100111101101011101001100001100110001011100001100101010111110100011010100111110000100000100111101000000010111001111101110010010111100111110000010011101001001000111011000010101010001011",
42 => "010011101010011101011000000010100000100100100111110100001000110010001011011010011101010000101111000111010011001011011100010101011110010001110000101100110000001001010010001000001101101101011010000001000001110010001111000101100100110111100000111011110110011",
43 => "100000000111011101001110000000011000111110100001111100101011100110011000101100010010110000001101010010110110000010001101001011000010100101000010100010110111100011010010011000110001000010000011000111001011101111001101001011011101010110000000110001011010100",
44 => "111010001111100000110000101010101101011001010000000011011110010110001011001110110101111010000101011010110001010100100100010000001111000110010010000010011000111101101011100001011111100011011101011001010000011011111011011111110011111110000111100000000000011",
45 => "100110101010010010110010001001100001101000010111001010010000100001000000111111111001100101110101100111001011101101100010100101010001001101011001110101011111000001110100010010101100011011110110011011011110010100010110100001001111010100111101100111111010011",
46 => "001011110100011001110001001110011100011010100101011100010001001011001000110001101000110100100000000100101001100000001110011110111000100100100110011101011110011001110110011100001110010110110001111001101111010110111110010100100000111110110000011010101010111",
47 => "010001100011010001101011001000001111010110001101001001010111110000000100000010101101010110100001110000010100101101101111000110110111000001101111111010110110001111000010111001011101111010110111100010111101010011010011011001001111100100101111101110110000000",
48 => "111100011110110101101000100011000100110010011011100100111110001100111110111000101000110011011000101111011010001010001110111001100111100001011110100101101001010001011011001001101110111101001110110111111100011101111110110011011101010001010010010100011010011",
49 => "111001101001111110100100001110010111110000101000000010110110101110001000100001010100111111000111000011110110111010100000001100000000001110011000101110000011100010010110111011000110000000001111001010000000101110001010100100010000101001001110000101110111000",
50 => "001101000101001010001101111110101011010000000010001101110111010100010011010101101001110101010001100111111111101111111111000110010001101110110110101110101110000110001000111110101000011001101001001000111000110001000100111001111100011001111110110000000000101",
51 => "000011110011000011000000101100000111111011001111100100001000110111111010100101011101000010101011100111100011110110100111101011111101010000101010111010101000011000101110010110100100010110000110010000000011001010000010001110000100000101111010101100100010011",
52 => "100010010100011111101101010011011001100010110011001001110101101001000010101001000001000000011000100111000001110001000100101111101100101010001111000100110010110101101100011010011101111001111100001111101110100001110011110100101000101010001010010100111010010",
53 => "001101101010001111100011001010000101010000010101111010000101111111000111011110001011111011000100111010001100101100010001100010000100000101001111001010101111111101000011101100001101110000000010010110101001001100111111110010011001100110110110101011000100101",
54 => "111101111101110100100100101010000101001111001111111100000101010111100111110011011011000011000011000000011111111000001010011111011011101000101011011001001010010100101010101010011000100000010110100100011000111010101001101110010101100111111000101110000111111",
55 => "100100001000111111100001000000111111010001010010100010100011011101010001101001100111011100001111011001010001100111111000011011000110010010101111011101111001010011011000110010010100010000010010101101000101110111111011110110111100111011101000111001101011010",
56 => "010100000001101000110100010000111001000011010111001010010110110011000100000101111111111100110010001001001101011111111110000011010110001100011001101100010100000110010110010000111101000111110101001001100011111010100110101100111000101010010001001101000111111",
57 => "001010101001100000010011011100011010100001011000110001101100010101111100010100101110000101000100111001000110110010101111011101101110101100110111100001010001111010011001110011100111101000100000011000100111111011101001010000111111011111001000111000010100011",
58 => "110010010000111010110011000010100111110010000011110011001010001111011100111101011111100010110011100101111010110001101111000100000011010110010010000111110000101110001100011000100111011001010011010000101100010001011110000111100100101000111100010110101001110",
59 => "101011000110111101010011011100000011001101011000000100100111110100101110010000010011011111011011011011101000100100010101101000011111000100101100101110110101010001100111010110101001101010001100111011011000011110011111000101010011101010111000111011100100100",
60 => "000000101111010101011100100101001100111110101000101101011011111001101110110010100000100010100100110110110011100011011100001010011110100100010000010011110111100011001001110010110010011101110011001101101111111010110010100111011111011000001100100101101010100",
61 => "101110100000110011100010010000100010111001001110010101001111110001111110010101010101000010111000010001111111010110000100010111110011001100000110111010001010100111011011011011011101001011111101000101110001110111111100001001101000101111101010011000111111101",
62 => "000110111111000110111101011000110101101101010110111101000010101111011010101010001100000111110100101100001000010011100011001011100100000110100100010111101010110011001111000000001000101110111110101010001110110001011111111000111100000100100110100010001111101",
63 => "101111001100100101011100010100110011110001100000000000010000100001000101101011000110001000001001100101000110100111111001101110010110011000001001001010111111110101000010011001000111110100110110110001100101000000011000100001011010011110100110010100111100111",
64 => "100110100010001110010100011101000101111000100001110010110010111011011111110100110110010100101101010000000011101100111001011101000011101111010100010010001100011000001101100111011011100100111010101011010100100011101100111011110110100001000110000101110100010",
65 => "010001010001101001110101101000110001010010011101001001010001101001000101000010100010001001101101110100011010010110101001000011000111110111111101111010000011101101011011011101001001011101110010001001100000101010110111000010000001001010000101010011011001111",
66 => "111110100011001110000000110110001111010111010000010111101001100111010100100101011110001110010010000110010110100111100000100000011010001111010100111011101010000010111111011110111001000011010000001110110011010101111111001110111111010110101000010101110001110",
67 => "001101000101011010000010010101111111110001000100010100011010111001000110110011111110010011100011101111101100111010000011011010101110111011100000011101000000000110110011011000010011111100010110111010000100000101010111010101100001100110100101010101111010000",
68 => "110100010010000111000110001010001000001011010101010100000010111000110111010111111100110001000010101000110111100001100010101011011101000100101011001000111110011011110001001010111011001001011011001110010110111001111001111010000111100110100110110111010010000",
69 => "101011011100010101011101100101101100001010110110000011101010110010001010100110110101011100000111101101000111000001011001001100011111100000011100010010100111111100010101100001101001100101010011101111101111001010111001110000000110011110111111100101010110101",
70 => "110101001011111010111100101001011010001000100110010011001011100010011010010011000111001111111000101100111010110011000010111101000001001101100110110000001110101011110110101010111011010101100111011110000001100110100100101100011100110110111001001110101011001",
71 => "111101111101111110000011001010001110011011001100011000000110101001000001011011100110010011100010000000101001111111010101000111111100010100101010111111010100010010101101001101111100100000000000110000101000001110100001110110010100011110010010100000101101110",
72 => "011110011000001101010011000001110110011110111001110000101100001001000001100101011110001001101100110101100110100111001011111000000000000101100101011101010100100001010001001110101101001101000111010111010000010011001011100000111010110101101010100001011101111",
73 => "001100010110110010001110000011101000001101110000111010100011000110111011010101101101010101111111011000000000111111011101100010110100000001000110011100001100010010010010001010110011011111111100100001111101100111011001111000111100010000011001111010000111001",
74 => "010111000010011010001000011010110010000011110011000000110100100110011010011101110011011010001010011111000000101101010000010000011000001011010001010100110101110010011001101011110111011001011011110101000110011010011100100011000110101100001100110101111010100",
75 => "100100111011000010111001110011100110110000000011101010111100010010100101001010000010110011001100010110011100010100100101101010101101100001101111010010111111000001001110100001100001000001000100001101101100010000111110000001001111100111110001000111101111011",
76 => "010110001010101010001110101001110101011101111110111111011110100000110011001011100011111011111000010111000111111100011000101001101000111000010110111101001111100011100110011001101001010011110010001101101010000110011110101111101101111111111000000011110100110",
77 => "111100100011000100111011011010001100011111111110011010111000000000010001001000110011001111010101110010111001001011101100111110110111001010011001111111010010000011001000011000011111010000011001011101010000101101011000001011101101001101001011111101100011000",
78 => "011000000011110100010111001011100001100110010100100010111110111001110101000001111110001001001000000011010111100010100011111101101110001110000110110100100001010001011101111011111111110110001111010111100101111010111001010010100110101001100001101111011111100",
79 => "110001000011110100101010010000011000010100111010001110010010001100000110101111010010101010000010001111110011110001011111010111011100111011111001001000111100011111010101101100000101011011100111111011011100110000011000011010101100101010111010100110110011100",
80 => "010110011100101100100011101100001101010100011011011101110001101101110100110100111011011110101110100110000110111100111001100100110101101011110110001110001100110111100110100000110010000011111111010101101110100010011000000110110111101110101001000010101101100",
81 => "001100001111100110010001111110100001100101011011010011110001010001011001100101010111011110011100110011000010000100011110111100010100100100011100111001101100010111100010001010000001000000011111111010101111110100011101100011001010101100011001000000000010001",
82 => "101011010100101100101100010101110110100111111010010000110111100000010110110110011101000011110000100011010001101110100000001010101111101110111110101001011011000011010000000101101101110110010001110111011010000000111101001111011100000010110100010011010010011",
83 => "110011111001101011010011001000100011000110010100011000101011110101000110100011101110000010010101010101001111111000100011000000000111010000001010111111111110101100011100110011110011001110111110011010111100001100011011100101110001011000111111000000011111101",
84 => "110000110011101110100001100001000110001110110101011001011010001101111110010101010111011100100110101001110101111000101010100001011110111101101011100101001010001110001110001011011110011010111011010010000101110001101010101001001010100110011101101110010100110",
85 => "011001101010011100000111011011000010011100000010010001100001011111101011110000100011101011110101001001100000100001001001001100110110001011110011101000111100010010111100010001010111001100111011111010100101001111010111001101111100011011001001100001110010100",
86 => "100101011101100110101111011111001000101011011111011001110100110001111011001101101101111010101000000110000001001100010100110001101110000011101110101001000101101100011011001100101111000101100000110001001000101011001010110001110010110111100110010010101010111",
87 => "100100000100001111100000000100100110000100110110010111011000000011000100011000100010010111100010011000101100110100101000011011011100101110001100011011011110010100011111100001010001100101011101011000111001001001110000001100001001101000110100011110010011001",
88 => "001110100100011001010010101111101101010101110001000101000101011000111000110000111110110110010111010010100010111111001000100010101000011111101110111101100111011110011111100011100001101011100100100000110100001011011000110100000110101001101111110010011000110",
89 => "101010010110101010011010001111100010011000001100100010101000100010011000111011110111011110010011100000100101000100000010101010101001000010000110100010101100011010001011100001100001110010010111101010111011001111100010101101101100110011010101101011001110110",
90 => "001001100011000110001000111111000001101001011101011001000101011111111111010011111011000001100011010110010111101001010011111000100110011101001111001111000110000001101001100010001000011010110010101011011111100100100100111011010101110000111010100100100100010",
91 => "101101101100100011111101100101001100000100001100110100110101000110011110100101100011000111111000110010111111111100110011010010001101011101000111010000010110111011110001010101011011100011111110011110000101101101100101010001110010110011100110011000000110110",
92 => "011111001100000111000110111110011011111001100100111110001100010001000100000001110110110111011001000011001011110001101100111101110100100100010011010000111001110001011000011110011100100110110011011101101010110010100111010001000101101011001110000001011110100",
93 => "010000011000011010100111000011101001000010110011100111011001100001001011111000110111100011101100001010100001010110001000000010111010010100110101000110001111100110010101000000101010010000101111101000011010010100001010110110101110000001010100011111010000010",
94 => "001100010100010100011100111000100110010011110110010111101000110111111100100110011100011101100000111110010001110100010100100110111110000101100011011110001110010111010001000101110100110001011011101111010111111101110110001100010110110011010100001000000110110",
95 => "111111011101111000001000000111100110110001010101101110000000111001101110001010011001001000000111100010011100000111100011001110101111100010000001111100011010100010001001101000011110010001100100101000110001011100100000001000100110110111100110110010101100100",
96 => "101111110000111110000000100001101101111111010110000110011010000011011101101111001011000010111110000010100101010111001101011101101001111101010111111010001101101101101101010000110111011110101011100100001000010100000111100000001011111110110011111010011001001",
97 => "111100101000001001010110011010000000000101101101101010111100101010110000111010010010011001111000001001000110110001111101010011001000010001011100101111011010111101001100110000101101101110100010101110111100010110001101001000111101110100010001111111000110101",
98 => "110011100111110111010101110100111001011011111011101000111011101001000100011000111101000100101001111111001001100000000011010110111010101001110111101100101001011100110101100010101101110001110011011010110011100011100111101000001000100000100010100010011000101",
99 => "001100010101010000000011111111110101010010110000110110001100010100100111100011000111011000100001010011100011010110011001011000110110101001100011000111000010001101001100111110111110110101110111011000101110001011111001001010110011010101001111111010110101011",
100 => "010100010100001111101010101011100001110101000101010011000111011010101011110100001000010111111111100011101111101110010010010011111111100101001110011110011101010000111001010000101001010011111101111001110111001100000111001111101110110000100101010001111000100"
);


constant ROM_R : ROM_type := ( 1 => "101101101000001000101000000101101000010001011010110010000100001000110101111011110000000101010001000011101010101011101000100111111000100101000100000110110000000110110010110110110100000000010011001001000010001010011000010011110100001110001011001100101111101",
2 => "010011111110111100101000101011111010001101110000110001000001111100010011111000000100011111101110000010001010110111011000110010111001111110110000111011101101100001011101111110110011001000011010111101100100110110001011100010100101100000110101011101011011010",
3 => "010000000110100101111010010000000011001100010110101000110110011011010111100001110111011100001110001010010001000001000000011000011001101011001000000001101111111000010010101001100110011100011110010001110110011101101001111000110000101110001111111000110111110",
4 => "011010011111001010111000110100001110100011110000001100001111101010001101001110111110100111111000111001111100110000010011000110111110010111111001000000100100010111111000010010001010101001100001110101111010111111101000101011101111010111101000010110110111101",
5 => "101101000010000110010110000000110001001000110101010110101000100110111100111011010110101100100111011000100100111111100010111110110111100110001011001101000001100011110000100101011001010101000011000000110110001101101000000011111000010101111010110111110110101",
6 => "001000100001110110011110101100110001110101110010000101010011100110111010110001000111001011100001101010011101101000111000001001111111000010100000000111000111111000111011101100101010111000111110100111111101101010100010100001000000000110010000110100011011101",
7 => "101111010010101010111010110111100111001111001111010101011101100011001101100101000111011101000011111000110100010001000011010010110101010100010111000110000111010010101001101010110001010000000010000101010010100101000011010010110100000110100010000101011000011",
8 => "010000111001000100000101011101110110001011101111110000010011110111110100011110001010010000111000111110101100000101011000100000101100111001000111110100110010101100001010101101101101000001000101100000010000101100101000001011011001011001101101011110110000010",
9 => "101000011100000101011111000001001011011010010110100001011101101001010101011011110010101001001101101001111001001110100000001100101100111100011111101111111100011000101110111100011100000011011001000111010100010111111100000001100011001110010000010001100111001",
10 => "100110111110101101001111011011000110000000101011011001000000100100111111001000101010011101100011010111101000000111111101101100011010101001111000000001010110010101010101111011111001101000111010100111111100101100101011101011101111101111111110111001001111101",
11 => "110010101001001000100100110001110001011110001111100011000010100100010100000000110110011001101001100011111010000111011100011011101111111000111001001100011110010001100111100000001100111001000001000000011110110011100010100010000101111010101010101010001000000",
12 => "110010000001110001001010101011100001110111111010111010101011111110010100010101111001011011010011011000111010110001110011100011001001000000110110000110011101110100000001001000101100011001011100010000111001101111111111110101011100001111011110111010011100001",
13 => "011011000110100011101011100000000111000000100010010001110010100000010110000001101101101101011111010110001000100110110110011011010101110110011111110000101110001101110001011011011101110100010110010010000110100011000011100110011001111101001100111001101011111",
14 => "010101101001110010101000011101110011110011111100010100011001010010101101111011001100010100100110010101111000110000001001100100000101110010101001111001011111100011010111111111100100111001001101100110110000000000001011011110000001100101000000010101111111100",
15 => "110100011111100011001111101111001001000001111100111101110110100111001011001001011000000001000111011100111011100100000000111100101001000011000001101100111101011100010000101010111001001100111001110000101110010100010000010111101001111000101100101100000010001",
16 => "110011100000001010110000100000000011100010011111001111101110100101111111101001110101000000011101111101000000100011010100111110111110101010000001000111111010001100111000010100010100010001101000101000111011110001111110001000101011001111111001101111010010111",
17 => "110000010111011100001111100000001001111100000111111000011011110101101111111100011100100010100100010101101110010101001010110011011000111101101111000110100111101010110111100000001101011111110000110101001111000001000011110011111110101111001010000001010001000",
18 => "010110100000110011010111101000010001100101001111100010110000010110100001010110000110001111011111001000110000111101110011100111101110111001001100000011001101001111101000000000110111111110101000011011000111011000011000101110111000101001111111100111010000011",
19 => "001010000100001110111011110101101101000000101001100010110010101000000011011000001111100110100101010100111100000100010111101100111000101010011111111111111010010000011001100011001010000011100101000100110111101100010011111001000010111000110100110000000011111",
20 => "000010110101101000111110100001000011001000111010000111111010100011011110110100001010110001001001010111110111100100101001001100111010001010110011001010011111000000101010111101000001110010100000111010100111110100101101011000101011001010000001000111111101111",
21 => "010000101000100101110100111011001001011100110000011010000100110011001001001111011100111011010110000010010010100000010101000111100010001001011111010010100100011011101110110100101110000001110100111110001001011001011101110011010010011000110011100000001010001",
22 => "011100001000111111011101010111111100010110110010111001011011101101111011001101000101001011101111001110011010101011010111111110001010010100000110001011011011111110010010100111011010011100011001011001101001110010010101011001100111101101001110100000011100011",
23 => "111111101100110101001101001010010000010011100101100100110100101100000010011111100100110111101001111100000101100011010101111101110110011110000010010101001000100110011111011001010000001001111110101100001010000100001110100111100001101000010110000110010100100",
24 => "100011110110111110011001101010011011110100010111111001011011000110010111101010100001111100111100111000001100100110101001001010101101100000101110000111010101111001001010101010111000101010001111110011101001100010111100110010011110010101100001110110001110100",
25 => "011101001010100111110001100001111110100010010011101001010101010100010011010001111001001010110100011011110101010101011100010001000011101000110111010001000101111001000000001011100101000110000101010111001111101001110101101011001101000110000010011100110010110",
26 => "100010100101001000001001010100011100001111001010111001011000110101111101000010001111010101110000011100111110001111111001001000101111111110010100100001111010010001001001110101110110101100111011101100111110000100101011110111011100111101000010000111111101010",
27 => "100001011110000010100010111110100110011101111100001101110101100101101001000101101101001101010101110111001111011101001110110010101101100100010011100111010000010000000101100110000101111011010101111000010110001111000000100000000010000101111111010011001010011",
28 => "010011011010001100010110011110101011100000101011100100111110010000111011110111001011001010101110111011011100101111010011101011011110010111100000110100000000110100100001111101011100100001111110101011011100000001000000101001001111110010100011101001101010111",
29 => "000110100101110011111110011110110010111001111111100110101100010100000010010101100110101110011011110110011011100111101101111000000100001111000011101111000010110101110000000010000101000011100101000010000100100001011101100000010000101001101011011100111011110",
30 => "011010100110101010100010011101101000000110101111100001000111111001001011011011011001110101110100101001011110101000001110101101001111100111111000010101001001010110011000000000001011001100101010011010010001101000100000100110101111110101100100101010100101001",
31 => "101111111110100100011010000011000101100001001101100110100101000011001000101100111010100000001111001010100101010110001100000000001000011001100110111010100001111001001010010010111110000110111001010011001000001000011110100010100010000010101111000110110001100",
32 => "010101101001011101010100001010111010100001100000000001001101100100111111100001011011000111001000111011111001101010001111001000000110101000100000010010111101101011000011001101001001001001001101000111010101110101001000110110110110111010000011110101111100001",
33 => "110100011011000010100011110111001000000010000010110110011100000110111000001000101000001010011001001100011010110010100101010100001101000101011000100101010011010110111110000101001100001100011010000100110100100010000101000101100100101011110100010101110000001",
34 => "010011111000001010001001000110111011111110110010000001110011111110100000010010101001011000110001111100010001000110001011100001111110100111010110010100101101001100111000101111111001001110101001110110001110111110100111110011100011111000101000010110100101000",
35 => "100111110111001110000000011111101010000111110100001000011111110100100000100111000001100110110000011011010001101111011011101000101011101010100100111001010111000110100001000011111011101000100101000000010100000111101001000001001000110111101110110011001101111",
36 => "000000001000101011101001111101001011101000110000000110110101101100110010001011101001111000000110111110101010110100100011111010010101000101010010001101110101111111110111110100001000000010010001010000111110000100010110000101111111000001100000101001001010100",
37 => "001100100101111110111010011010011010110011000010011001000100011100001111001001110110100101011100000000110111001101101101101110100011100010001101111101011011010001100100000111010010110010101010011101010011011000010111100010010101100001100110101011010001010",
38 => "111010011110011010101001101010011001100000111001100100111010100010001011110000001010010100111111111000111010001100011110000111101011100100010000000101000110011100010011010110111111001000101111011111101011001100110011001101100000011101011011001111001001111",
39 => "100000011110010101010110100001010110011011100011010011010110100001010001011101110100010010010111100111110101010101011010010111001101111001000110101100100110000001000101010011010010010111010101010011011001111100001011101001100100110111001010010000000000000",
40 => "111100100111001001000000011101011010000111110010000101001011100110110101111100111000100101101001010110000111110001110000000100001001010110100101000100110010101110100010000000000000101011101101111110101001001111000010101011110111011001010001111000100011001",
41 => "001101110101010100001011000100001101100101111101011000001010111110001101100111101101011101001100001100110001011100001100101010111110100011010100111110000100000100101101000000010111001111101110010010111100111110000010011101001001000111011000010101010001011",
42 => "010011101010011101011000000010100000100100100111110100001000110010001011011010011101010000101111000111010011001011011100010101011110010001110000101100110000001001010010001000001101101101011010001001000001110011001111000101100100110111100000111011110110011",
43 => "100000000111011101001110000000011000111110100001111100101011100110011000101100010010010000001101010010110110000010001101001011000010100101000010100010110111100011010010011000110001000010000011000111001011101111001101001011011101010110000000010001011010100",
44 => "111010001111100000010000101010101101011001010000000011011110010110001011001110110101111011000101011010110001010100100100010000001111000110010010000010011000111101101011100001011111100011011101011001010000011011111011011111110011111110000111100000000000011",
45 => "100110101010010010110010001001100001101000010111101010010000100001000000111111111001100101110101100111001011100101100010100101010001001101011001110101011111000001110100010010101100011011110110011011011110010100010110100001001111010100111101100111111010011",
46 => "000011110100011001110001001100011100011010100101011100010001001011001000110001101000110100100000000100101001100000001110011110111000100100100110011101011110011001110110011100001110010110110001111001101111010110111110010100100000111110110000011010101010111",
47 => "000001100011010001101011001000001111010110001101001001010111110000000100000010101101010110100001110000010100101101101111000110110111000001101111111010110110001111000010111001011101111010110111100010111101010011010011011001001011100100101111101110110000000",
48 => "111100011110110101101000100011000100110010011011100100111110001100111110111000101000110011011000101111011010001010001110111001100111100001011110100101101101010001010011001001101110111101001110110111111100011101111110110011011101010001010010010100011010011",
49 => "101001101001111110100100001110010111110000101000000010110110101110001000100001010100111111000111000011110110111010100000001100000000001010011000101110000011100010010110111011000110000000001111001010000000101110001010100100010000101001001110000101110111000",
50 => "001101000101001010001101111110101011010000000010001101110111010100010011010101101001110101010001100111111111101111011111000110010001101110110110101110101110000110001000111110101000011001101001001000111000110001000100111001111100011001111110010000000000101",
51 => "000011110011100011000000101100000111111011001111100101001000110111111010100101011101000010101011100111100011110110100111101011111101010000101010111010101000011000101110010110100100010110000110010000000011001010000010001110000100000101111010101100100010011",
52 => "100010010100011111101101010011011001100010110011001001110101101001000010101001000001000000011000000111000001110001000100101111101100101010001111000100110010110101101100011010011101111001111100001111001110100001110011110100101000101010001010010100111010010",
53 => "001101101010001111100011001010000101010000010101111010000101111111000111011110001011111011000100101010001100101100010001100010000100000101001111001010101111111101000011101100001101110000000010010110101001001100111111110010011001000110110110101011000100101",
54 => "111101111101110100100100101010000101001111001111111100000101010111100111110011011011000011000011000000011101111000001010011111011011101000101011011001001010010101101010101010011000100000010110100100011000111010101001101110010101100111111000101110000111111",
55 => "100100000000111111100001000000111111010001010010100010100011011101010001101001100111011100001111011001010001100111111000011011000110010010101111010101111001010011011000110010010100010000010010101101000101110111111011110110111100111011101000111001101011010",
56 => "010100000001101000110100010000111001000011010111001010010110110011000100000101111111111100110010001001001101011111111110000011010110001100011001101100010100000110010110010000111101000110110101001001100011111010101110101100111000101010010001001101000111111",
57 => "001010101001100000010011011100011010100001011000110001101100010101111100010100101110000101000100111001000110110010101110011101101110101100110111100001010001111010011001110011100111001000100000011000100111111011101001010000111111011111001000111000010100011",
58 => "110010010000111010110011000010100111110010000011110011001010001111011100111101011111100010110011100101111010110001101111000100000011010110110010000111110000101110001100011000100111011001010011010000101100010001011110000111100100101000111100000110101001110",
59 => "101011100110111101010011011100000011001101011000000100100111110100101110010000010011011111011011011011101000100100010101101000011111000100101100101110110101010001100111010110101001101010001100111001011000011110011111000101010011101010111000111011100100100",
60 => "000000101111010101011100100101001100111110101010101101011011111001101110110010100000100010100101110110110011100011011100001010011110100100010000010011110111100011001001110010110010011101110011001101101111111010110010100111011111011000001100100101101010100",
61 => "101110100000110011100010010000100010111001001010010101001111110001111110010101010101000010111000010001111111010110000100010111110011001100000110111010001010100111011011011011011101001011111101000101110001110111111100000001101000101111101010011000111111101",
62 => "000110111111000110111101011000110101101101010110111101000010101111011010101010101100000111110100101100001000010011100001001011100100000110100100010111101010110011001111000000001000101110111110101010001110110001011111111000111100000100100110100010001111101",
63 => "101111001100100101011100010100110011110001100000000000010000100001000101101011000110001000001001101101000110100111111001101110010110011000001001001010111111110101000010011001000111110100110110110001100101000000011000100001011010011110100110011100111100111",
64 => "100110100010001110010100011101000101111000100001110010110010111011011110100100110110010100101101010000000011101100111001011101000011101111010100010010001100011000001101100111011011100100111010101011010100100011101100111011110110100001000110000101110100010",
65 => "010001010001101001110101101000110001010010010101001001010001101001000101000010100010001000101101110100011010010110101001000011000111110111111101111010000011101101011011011101001001011101110010001001100000101010110111000010000001001010000101010011011001111",
66 => "111110100011001110000000110110001111010111010000010111101001100011010100100101011110001110010010000110010110100111100000100000011010001111010100111011101011000010111111011110111001000011010000001110110011010101111111001110111111010110101000010101110001110",
67 => "001101001101011010000010010101111111110001000100010100011010111001000110110011111110010011100011101111101100111010000011011010101110111011100000011101000000000110110011011100010011111100010110111010000100000101010111010101100001100110100101010101111010000",
68 => "110100010010000111000110001010001000001011010101010100000010111000010111010111111100110001000010101000110111100001100010101011011101000100101011001000111110011011110001001010111011001001011011001110010110111001111001111010000111100110100110110111010010010",
69 => "101011011100010101011101100101101100001010110110000011101010110010011010100110110101011100000111101101000111000001011001001100011110100000011100010010100111111100010101100001101001100101010011101111101111001010111001110000000110011110111111100101010110101",
70 => "110101001011111010111100101001011010001000100110010011001011100010011010010011000111001111111000101100111010110011000010111101000001000101100110110000001110101011110110101010011011010101100111011110000001100110100100101100011100110110111001001110101011001",
71 => "111101111101111110000011001010001110011011001100011000000110101001000001010011100110010011000010000000101001111111010101000111111100010100101010111111010100010010101101001101111100100000000000110000101000001110100001110110010100011110010010100000101101110",
72 => "011110011000001101010011010001110110011110111001110000101100001001000001100101011110001001101100110101100110100111001011111000000000001101100101011101010100100001010001001110101101001101000111010111010000010011001011100000111010110101101010100001011101111",
73 => "001110010110110010001110000011101000001101110000111010100011000110111011010101100101010101111111011000000000111111011101100010110100000001000110011100001100010010010010001010110011011111111100100001111101100111011001111000111100010000011001111010000111001",
74 => "010111000010011010001000011010110010000011110011000000110100100110011010011101110011011010001010011111000000101101010000010000011001001011010001010100110101110010011001101011110111011001011011110101000110011010011100100011000110101100001100110101111010101",
75 => "100100111011000010111001110011100110110000000011101010111100010010100101001010000010110011001100010110011100010000100101101010101101100001101111010010111111000001001110100001100001000001000100001101101100010000111110000000001111100111110001000111101111011",
76 => "010110001010101010001110101001110101011101111110111111011110100000110011001011100011111011111000010111000111111100011000101001101000111000010110111101001111100011100110011001100001010011110010001101101011000110011110101111101101111111111000000011110100110",
77 => "111100100011000100111011011010001100011111111110011010111000000000010001001000110011001111011101110010111001001011101100111110110111001010011001111111010010000011001000011000011101010000011001011101010000101101011000001011101101001101001011111101100011000",
78 => "011000000010110100010111001011100001100110010100100010111110111001110101000001111110001001001000000011010111100010100011111101101110001110000110110100100001010001011101111011111011110110001111010111100101111010111001010010100110101001100001101111011111100",
79 => "110001000011110100101010010000011000110100111010001110010010001100000110101111010010101010000010001111110011110001011111010111011100111011111001001000111100011111010101101100000101011011100111111011011100110000011000011010001100101010111010100110110011100",
80 => "010110011100101100100011101100001101010100011011011101110001101101110100110100111011011110101110100110000110111100111001100100110101101011110110001110001100110111100110100000110010000011111111010101101110100110011000000110110111101111101001000010101101100",
81 => "001100001111100110010001111110100001100101011011010011110001010001011001100101010111011110011100110011100010000100011110111100000100100100011100111001101100010111100010001010000001000000011111111010101111110100011101100011001010101100011001000000000010001",
82 => "101011010100101100101100010101110110100111111010010000110111100001010110110110011101000011110000100011010001101110100000001010101111101110111110101001010011000011010000000101101101110110010001110111011010000000111101001111011100000010110100010011010010011",
83 => "110011111001101011010011001000100011000110010100011000101011110101000110100011101110000010010101010101001111111000100011000000000111010000001010111111111110101100011100110011110011001110111110111010111100001100011011100101110001011000111111000000111111101",
84 => "110000110011101110100001100001000110001110110101011001011010001101111110010101010111011100100110101001110001111000101010100001011110111101101011100101001010001110001110001011011110011010111011010010000111110001101010101001001010100110011101101110010100110",
85 => "011001101010011100000111011011000010011100000010010001100001011111101011110000100011101011110101001101100000100001001001001100110110001011110011101000111100010010111100010001010111001000111011111010100101001111010111001101111100011011001001100001110010100",
86 => "100101010101100110101111011111001000101011011111011001110100110001111011001101101101111010101000000110000001001100010100110001101110000011101110101001000101101100011011001100101111000101100000110001001000101011001010110001110000110111100110010010101010111",
87 => "100100000100001111100000000100100110000100110110010111011000000011000100011000100010000111100010011000101100110100101000011011011100101110001100011011011110010100011111100001010001100101001101011000111001001001110000001100001001101000110100011110010011001",
88 => "001110100101011001010010101111101101010101110001000101000101011000111000110000111110110110010111010010100010111111001000100010101000011111101110111101100111011110011111100011100001101011100100100000110100011011011000110100000110101001101111110010011000110",
89 => "101010010110101010011010001111100010011000001110100010101000100010011000111011110111011110010011100000100101000100000010101010101001100010000110100010101100011010001011100001100001110010010111101010111011001111100010101101101100110011010101101011001110110",
90 => "001001100011000110001000111111000001101001011101011001000101011111111111010011111011000001100011010110000111101001010011111000100110011101001111001111000110000001101001100110001000011010110010101011011111100100100100111011010101110000111010100100100100010",
91 => "101101101100100011111101100101001100000100011100110100110101000110011110100101100011000111111000110010111111111100110011010010001101011101000111010000010111111011110001010101011011100011111110011110000101101101100101010001110010110011100110011000000110110",
92 => "011111001100000111000110111110011011111001100100110110001100010001000100000001110110110111011001000011001011110001101100111101110100100100010011010000111001110001011000011110011000100110110011011101101010110010100111010001000101101011001110000001011110100",
93 => "010000011000011110100111000011111001000010110011100111011001100001001011111000110111100011101100001010100001010110001000000010111010010100110101000110001111100110010101000000101010010000101111101000011010010100001010110110101110000001010100011111010000010",
94 => "001100110100010100011100111000100110010011010110010111101000110111111100100110011100011101100000111110010001110100010100100110111110000101100011011110001110010111010001000101110100110001011011101111010111111101110110001100010110110011010100001000000110110",
95 => "111111011101111000001000000111100110110001010101101110000000111001101110001010011001001000000111100010011100000011100011001110101111100010000001111101011010100010001001101000011110010001100100101000110001011100100000001000100110110111100110110010101100100",
96 => "101111110000111110000000100001101001111111010110000110011010000011011101101111001011000010111110000010100101010111001101011101101001111101010111111010001101101101101101010000110111011110101011100100001001010100000111100000001011111110110011111010011001001",
97 => "111100111000001001010110011010000000000101101101101010111100101010110000111010010010011001111000001001000110110101111101010011001000010001011100101111011010111101001100110000101101101110100010101110111100010110001101001000111101110100010001111111000110101",
98 => "110011100111110111010101110100111001011111111011101000111011101001000100011000111101000100101001111111001001100000000011010110111010101001110111101100101001011110110101100010101101110001110011011010110011100011100111101000001000100000100010100010011000101",
99 => "001100010101010000000011111111110101010010110000110110000100010100100111100011000111011000100001010011100011010110011001011000110110101001100011000111000010001101001100110110111110110101110111011000101110001011111001001010110011010101001111111010110101011",
100 => "010100010100001111101010101011100001110101000101010011000111011010101011100100001000010111111111100011101111101110010010010011111111100101001110011110011101010000111001010000101001010001111101111001110111001100000111001111101110110000100101010001111000100"
);


begin

CLOCK_PROGRESS : process
	begin
		Clock<='0';
		wait for clk_period/2;
		Clock<='1';
		wait for clk_period/2;
end process;

tester : process (Clock)
begin

	--test <= ROM_R(0);
	--check <= ROM_C(0);

	if (counter = 100) then
		counter <= 1;
		test <= ROM_R(counter);
		check <= ROM_C(counter);
	else
		counter <= counter + 1;
		test <= ROM_R(counter);
		check <= ROM_C(counter);
	end if;

end process;


checker : process (Clock,result)
begin
	if (result = check) then
		ok <= '1';
	else
		ok <= '0';
	end if;
end process;


dut : Decoder
	port map(
		clock  => Clock,
		input	=> test, --ROM_SINGLEin(0), --test,
		output => result
	);

end architecture;