--mads
LIBRARY IEEE;
USE IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.std_logic_unsigned.all;

entity DecoderBCHEModSumHelper is
	port(  
		input  : in std_logic_vector(254 downto 0);
		output : out std_logic
	);
end entity;

architecture DecoderBCHEModSumHelper_arch of DecoderBCHEModSumHelper is

type ROM_typeMOD is array (0 to 255) of integer;
constant ROM_MOD2 : ROM_typeMOD := ( 0 => 0,
1 => 1,
2 => 0,
3 => 1,
4 => 0,
5 => 1,
6 => 0,
7 => 1,
8 => 0,
9 => 1,
10 => 0,
11 => 1,
12 => 0,
13 => 1,
14 => 0,
15 => 1,
16 => 0,
17 => 1,
18 => 0,
19 => 1,
20 => 0,
21 => 1,
22 => 0,
23 => 1,
24 => 0,
25 => 1,
26 => 0,
27 => 1,
28 => 0,
29 => 1,
30 => 0,
31 => 1,
32 => 0,
33 => 1,
34 => 0,
35 => 1,
36 => 0,
37 => 1,
38 => 0,
39 => 1,
40 => 0,
41 => 1,
42 => 0,
43 => 1,
44 => 0,
45 => 1,
46 => 0,
47 => 1,
48 => 0,
49 => 1,
50 => 0,
51 => 1,
52 => 0,
53 => 1,
54 => 0,
55 => 1,
56 => 0,
57 => 1,
58 => 0,
59 => 1,
60 => 0,
61 => 1,
62 => 0,
63 => 1,
64 => 0,
65 => 1,
66 => 0,
67 => 1,
68 => 0,
69 => 1,
70 => 0,
71 => 1,
72 => 0,
73 => 1,
74 => 0,
75 => 1,
76 => 0,
77 => 1,
78 => 0,
79 => 1,
80 => 0,
81 => 1,
82 => 0,
83 => 1,
84 => 0,
85 => 1,
86 => 0,
87 => 1,
88 => 0,
89 => 1,
90 => 0,
91 => 1,
92 => 0,
93 => 1,
94 => 0,
95 => 1,
96 => 0,
97 => 1,
98 => 0,
99 => 1,
100 => 0,
101 => 1,
102 => 0,
103 => 1,
104 => 0,
105 => 1,
106 => 0,
107 => 1,
108 => 0,
109 => 1,
110 => 0,
111 => 1,
112 => 0,
113 => 1,
114 => 0,
115 => 1,
116 => 0,
117 => 1,
118 => 0,
119 => 1,
120 => 0,
121 => 1,
122 => 0,
123 => 1,
124 => 0,
125 => 1,
126 => 0,
127 => 1,
128 => 0,
129 => 1,
130 => 0,
131 => 1,
132 => 0,
133 => 1,
134 => 0,
135 => 1,
136 => 0,
137 => 1,
138 => 0,
139 => 1,
140 => 0,
141 => 1,
142 => 0,
143 => 1,
144 => 0,
145 => 1,
146 => 0,
147 => 1,
148 => 0,
149 => 1,
150 => 0,
151 => 1,
152 => 0,
153 => 1,
154 => 0,
155 => 1,
156 => 0,
157 => 1,
158 => 0,
159 => 1,
160 => 0,
161 => 1,
162 => 0,
163 => 1,
164 => 0,
165 => 1,
166 => 0,
167 => 1,
168 => 0,
169 => 1,
170 => 0,
171 => 1,
172 => 0,
173 => 1,
174 => 0,
175 => 1,
176 => 0,
177 => 1,
178 => 0,
179 => 1,
180 => 0,
181 => 1,
182 => 0,
183 => 1,
184 => 0,
185 => 1,
186 => 0,
187 => 1,
188 => 0,
189 => 1,
190 => 0,
191 => 1,
192 => 0,
193 => 1,
194 => 0,
195 => 1,
196 => 0,
197 => 1,
198 => 0,
199 => 1,
200 => 0,
201 => 1,
202 => 0,
203 => 1,
204 => 0,
205 => 1,
206 => 0,
207 => 1,
208 => 0,
209 => 1,
210 => 0,
211 => 1,
212 => 0,
213 => 1,
214 => 0,
215 => 1,
216 => 0,
217 => 1,
218 => 0,
219 => 1,
220 => 0,
221 => 1,
222 => 0,
223 => 1,
224 => 0,
225 => 1,
226 => 0,
227 => 1,
228 => 0,
229 => 1,
230 => 0,
231 => 1,
232 => 0,
233 => 1,
234 => 0,
235 => 1,
236 => 0,
237 => 1,
238 => 0,
239 => 1,
240 => 0,
241 => 1,
242 => 0,
243 => 1,
244 => 0,
245 => 1,
246 => 0,
247 => 1,
248 => 0,
249 => 1,
250 => 0,
251 => 1,
252 => 0,
253 => 1,
254 => 0,
255 => 1
);

type ROM_typeSum is array (0 to 255) of integer range 0 to 8;
constant ROM_SUM : ROM_typeSum := ( 0 => 0,
1 => 1,
2 => 1,
3 => 2,
4 => 1,
5 => 2,
6 => 2,
7 => 3,
8 => 1,
9 => 2,
10 => 2,
11 => 3,
12 => 2,
13 => 3,
14 => 3,
15 => 4,
16 => 1,
17 => 2,
18 => 2,
19 => 3,
20 => 2,
21 => 3,
22 => 3,
23 => 4,
24 => 2,
25 => 3,
26 => 3,
27 => 4,
28 => 3,
29 => 4,
30 => 4,
31 => 5,
32 => 1,
33 => 2,
34 => 2,
35 => 3,
36 => 2,
37 => 3,
38 => 3,
39 => 4,
40 => 2,
41 => 3,
42 => 3,
43 => 4,
44 => 3,
45 => 4,
46 => 4,
47 => 5,
48 => 2,
49 => 3,
50 => 3,
51 => 4,
52 => 3,
53 => 4,
54 => 4,
55 => 5,
56 => 3,
57 => 4,
58 => 4,
59 => 5,
60 => 4,
61 => 5,
62 => 5,
63 => 6,
64 => 1,
65 => 2,
66 => 2,
67 => 3,
68 => 2,
69 => 3,
70 => 3,
71 => 4,
72 => 2,
73 => 3,
74 => 3,
75 => 4,
76 => 3,
77 => 4,
78 => 4,
79 => 5,
80 => 2,
81 => 3,
82 => 3,
83 => 4,
84 => 3,
85 => 4,
86 => 4,
87 => 5,
88 => 3,
89 => 4,
90 => 4,
91 => 5,
92 => 4,
93 => 5,
94 => 5,
95 => 6,
96 => 2,
97 => 3,
98 => 3,
99 => 4,
100 => 3,
101 => 4,
102 => 4,
103 => 5,
104 => 3,
105 => 4,
106 => 4,
107 => 5,
108 => 4,
109 => 5,
110 => 5,
111 => 6,
112 => 3,
113 => 4,
114 => 4,
115 => 5,
116 => 4,
117 => 5,
118 => 5,
119 => 6,
120 => 4,
121 => 5,
122 => 5,
123 => 6,
124 => 5,
125 => 6,
126 => 6,
127 => 7,
128 => 1,
129 => 2,
130 => 2,
131 => 3,
132 => 2,
133 => 3,
134 => 3,
135 => 4,
136 => 2,
137 => 3,
138 => 3,
139 => 4,
140 => 3,
141 => 4,
142 => 4,
143 => 5,
144 => 2,
145 => 3,
146 => 3,
147 => 4,
148 => 3,
149 => 4,
150 => 4,
151 => 5,
152 => 3,
153 => 4,
154 => 4,
155 => 5,
156 => 4,
157 => 5,
158 => 5,
159 => 6,
160 => 2,
161 => 3,
162 => 3,
163 => 4,
164 => 3,
165 => 4,
166 => 4,
167 => 5,
168 => 3,
169 => 4,
170 => 4,
171 => 5,
172 => 4,
173 => 5,
174 => 5,
175 => 6,
176 => 3,
177 => 4,
178 => 4,
179 => 5,
180 => 4,
181 => 5,
182 => 5,
183 => 6,
184 => 4,
185 => 5,
186 => 5,
187 => 6,
188 => 5,
189 => 6,
190 => 6,
191 => 7,
192 => 2,
193 => 3,
194 => 3,
195 => 4,
196 => 3,
197 => 4,
198 => 4,
199 => 5,
200 => 3,
201 => 4,
202 => 4,
203 => 5,
204 => 4,
205 => 5,
206 => 5,
207 => 6,
208 => 3,
209 => 4,
210 => 4,
211 => 5,
212 => 4,
213 => 5,
214 => 5,
215 => 6,
216 => 4,
217 => 5,
218 => 5,
219 => 6,
220 => 5,
221 => 6,
222 => 6,
223 => 7,
224 => 3,
225 => 4,
226 => 4,
227 => 5,
228 => 4,
229 => 5,
230 => 5,
231 => 6,
232 => 4,
233 => 5,
234 => 5,
235 => 6,
236 => 5,
237 => 6,
238 => 6,
239 => 7,
240 => 4,
241 => 5,
242 => 5,
243 => 6,
244 => 5,
245 => 6,
246 => 6,
247 => 7,
248 => 5,
249 => 6,
250 => 6,
251 => 7,
252 => 6,
253 => 7,
254 => 7,
255 => 8
);

signal sum : integer range 0 to 255;
signal modsum : integer range 0 to 1;
signal test : std_logic_vector(255 downto 0);

begin

test <= "0" & input;

sum <= ROM_SUM(to_integer(unsigned(test(7 downto 0)))) +ROM_SUM(to_integer(unsigned(test(15 downto 8)))) +ROM_SUM(to_integer(unsigned(test(23 downto 16)))) +ROM_SUM(to_integer(unsigned(test(31 downto 24)))) +ROM_SUM(to_integer(unsigned(test(39 downto 32)))) +ROM_SUM(to_integer(unsigned(test(47 downto 40)))) +ROM_SUM(to_integer(unsigned(test(55 downto 48)))) +ROM_SUM(to_integer(unsigned(test(63 downto 56)))) +ROM_SUM(to_integer(unsigned(test(71 downto 64)))) +ROM_SUM(to_integer(unsigned(test(79 downto 72)))) +ROM_SUM(to_integer(unsigned(test(87 downto 80)))) +ROM_SUM(to_integer(unsigned(test(95 downto 88)))) +ROM_SUM(to_integer(unsigned(test(103 downto 96)))) +ROM_SUM(to_integer(unsigned(test(111 downto 104)))) +ROM_SUM(to_integer(unsigned(test(119 downto 112)))) +ROM_SUM(to_integer(unsigned(test(127 downto 120)))) +ROM_SUM(to_integer(unsigned(test(135 downto 128)))) +ROM_SUM(to_integer(unsigned(test(143 downto 136)))) +ROM_SUM(to_integer(unsigned(test(151 downto 144)))) +ROM_SUM(to_integer(unsigned(test(159 downto 152)))) +ROM_SUM(to_integer(unsigned(test(167 downto 160)))) +ROM_SUM(to_integer(unsigned(test(175 downto 168)))) +ROM_SUM(to_integer(unsigned(test(183 downto 176)))) +ROM_SUM(to_integer(unsigned(test(191 downto 184)))) +ROM_SUM(to_integer(unsigned(test(199 downto 192)))) +ROM_SUM(to_integer(unsigned(test(207 downto 200)))) +ROM_SUM(to_integer(unsigned(test(215 downto 208)))) +ROM_SUM(to_integer(unsigned(test(223 downto 216)))) +ROM_SUM(to_integer(unsigned(test(231 downto 224)))) +ROM_SUM(to_integer(unsigned(test(239 downto 232)))) +ROM_SUM(to_integer(unsigned(test(247 downto 240)))) +ROM_SUM(to_integer(unsigned(test(255 downto 248))));

process(sum)
begin
if (sum < 256) then
modsum <= ROM_MOD2(sum);
end if;
end process;

process(modsum)
begin

if (modsum = 1) then
	output <= '1';
else
	output <= '0';
end if;

end process;

end architecture;


